
module embedded_system (
	ad9833_io_readdata,
	clk_clk);	

	output	[31:0]	ad9833_io_readdata;
	input		clk_clk;
endmodule
