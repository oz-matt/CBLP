// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"

// DATE "01/12/2020 22:55:32"

// 
// Device: Altera EP4CGX150DF31C7 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module qtestpd (
	clk_clk,
	onchip_memory2_0_s1_address,
	onchip_memory2_0_s1_clken,
	onchip_memory2_0_s1_chipselect,
	onchip_memory2_0_s1_write,
	onchip_memory2_0_s1_readdata,
	onchip_memory2_0_s1_writedata,
	onchip_memory2_0_s1_byteenable,
	onchip_memory2_0_s2_address,
	onchip_memory2_0_s2_chipselect,
	onchip_memory2_0_s2_clken,
	onchip_memory2_0_s2_write,
	onchip_memory2_0_s2_readdata,
	onchip_memory2_0_s2_writedata,
	onchip_memory2_0_s2_byteenable,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
input 	clk_clk;
input 	[13:0] onchip_memory2_0_s1_address;
input 	onchip_memory2_0_s1_clken;
input 	onchip_memory2_0_s1_chipselect;
input 	onchip_memory2_0_s1_write;
output 	[63:0] onchip_memory2_0_s1_readdata;
input 	[63:0] onchip_memory2_0_s1_writedata;
input 	[7:0] onchip_memory2_0_s1_byteenable;
input 	[13:0] onchip_memory2_0_s2_address;
input 	onchip_memory2_0_s2_chipselect;
input 	onchip_memory2_0_s2_clken;
input 	onchip_memory2_0_s2_write;
output 	[63:0] onchip_memory2_0_s2_readdata;
input 	[63:0] onchip_memory2_0_s2_writedata;
input 	[7:0] onchip_memory2_0_s2_byteenable;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[0]~0_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[1]~1_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[2]~2_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[3]~3_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[4]~4_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[5]~5_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[6]~6_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[7]~7_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[8]~8_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[9]~9_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[10]~10_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[11]~11_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[12]~12_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[13]~13_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[14]~14_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[15]~15_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[16]~16_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[17]~17_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[18]~18_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[19]~19_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[20]~20_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[21]~21_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[22]~22_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[23]~23_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[24]~24_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[25]~25_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[26]~26_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[27]~27_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[28]~28_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[29]~29_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[30]~30_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[31]~31_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[32]~32_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[33]~33_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[34]~34_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[35]~35_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[36]~36_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[37]~37_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[38]~38_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[39]~39_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[40]~40_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[41]~41_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[42]~42_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[43]~43_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[44]~44_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[45]~45_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[46]~46_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[47]~47_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[48]~48_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[49]~49_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[50]~50_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[51]~51_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[52]~52_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[53]~53_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[54]~54_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[55]~55_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[56]~56_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[57]~57_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[58]~58_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[59]~59_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[60]~60_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[61]~61_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[62]~62_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[63]~63_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[0]~0_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[1]~1_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[2]~2_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[3]~3_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[4]~4_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[5]~5_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[6]~6_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[7]~7_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[8]~8_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[9]~9_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[10]~10_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[11]~11_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[12]~12_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[13]~13_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[14]~14_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[15]~15_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[16]~16_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[17]~17_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[18]~18_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[19]~19_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[20]~20_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[21]~21_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[22]~22_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[23]~23_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[24]~24_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[25]~25_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[26]~26_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[27]~27_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[28]~28_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[29]~29_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[30]~30_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[31]~31_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[32]~32_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[33]~33_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[34]~34_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[35]~35_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[36]~36_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[37]~37_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[38]~38_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[39]~39_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[40]~40_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[41]~41_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[42]~42_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[43]~43_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[44]~44_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[45]~45_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[46]~46_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[47]~47_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[48]~48_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[49]~49_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[50]~50_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[51]~51_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[52]~52_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[53]~53_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[54]~54_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[55]~55_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[56]~56_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[57]~57_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[58]~58_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[59]~59_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[60]~60_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[61]~61_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[62]~62_combout ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[63]~63_combout ;
wire \rst_controller|r_early_rst~q ;
wire \onchip_memory2_0_s1_address[13]~input_o ;
wire \onchip_memory2_0_s1_chipselect~input_o ;
wire \onchip_memory2_0_s1_write~input_o ;
wire \onchip_memory2_0_s2_address[13]~input_o ;
wire \onchip_memory2_0_s2_chipselect~input_o ;
wire \onchip_memory2_0_s2_write~input_o ;
wire \clk_clk~input_o ;
wire \onchip_memory2_0_s1_clken~input_o ;
wire \onchip_memory2_0_s2_clken~input_o ;
wire \onchip_memory2_0_s1_writedata[0]~input_o ;
wire \onchip_memory2_0_s1_address[0]~input_o ;
wire \onchip_memory2_0_s1_address[1]~input_o ;
wire \onchip_memory2_0_s1_address[2]~input_o ;
wire \onchip_memory2_0_s1_address[3]~input_o ;
wire \onchip_memory2_0_s1_address[4]~input_o ;
wire \onchip_memory2_0_s1_address[5]~input_o ;
wire \onchip_memory2_0_s1_address[6]~input_o ;
wire \onchip_memory2_0_s1_address[7]~input_o ;
wire \onchip_memory2_0_s1_address[8]~input_o ;
wire \onchip_memory2_0_s1_address[9]~input_o ;
wire \onchip_memory2_0_s1_address[10]~input_o ;
wire \onchip_memory2_0_s1_address[11]~input_o ;
wire \onchip_memory2_0_s1_address[12]~input_o ;
wire \onchip_memory2_0_s1_byteenable[0]~input_o ;
wire \onchip_memory2_0_s2_writedata[0]~input_o ;
wire \onchip_memory2_0_s2_address[0]~input_o ;
wire \onchip_memory2_0_s2_address[1]~input_o ;
wire \onchip_memory2_0_s2_address[2]~input_o ;
wire \onchip_memory2_0_s2_address[3]~input_o ;
wire \onchip_memory2_0_s2_address[4]~input_o ;
wire \onchip_memory2_0_s2_address[5]~input_o ;
wire \onchip_memory2_0_s2_address[6]~input_o ;
wire \onchip_memory2_0_s2_address[7]~input_o ;
wire \onchip_memory2_0_s2_address[8]~input_o ;
wire \onchip_memory2_0_s2_address[9]~input_o ;
wire \onchip_memory2_0_s2_address[10]~input_o ;
wire \onchip_memory2_0_s2_address[11]~input_o ;
wire \onchip_memory2_0_s2_address[12]~input_o ;
wire \onchip_memory2_0_s2_byteenable[0]~input_o ;
wire \onchip_memory2_0_s1_writedata[1]~input_o ;
wire \onchip_memory2_0_s2_writedata[1]~input_o ;
wire \onchip_memory2_0_s1_writedata[2]~input_o ;
wire \onchip_memory2_0_s2_writedata[2]~input_o ;
wire \onchip_memory2_0_s1_writedata[3]~input_o ;
wire \onchip_memory2_0_s2_writedata[3]~input_o ;
wire \onchip_memory2_0_s1_writedata[4]~input_o ;
wire \onchip_memory2_0_s2_writedata[4]~input_o ;
wire \onchip_memory2_0_s1_writedata[5]~input_o ;
wire \onchip_memory2_0_s2_writedata[5]~input_o ;
wire \onchip_memory2_0_s1_writedata[6]~input_o ;
wire \onchip_memory2_0_s2_writedata[6]~input_o ;
wire \onchip_memory2_0_s1_writedata[7]~input_o ;
wire \onchip_memory2_0_s2_writedata[7]~input_o ;
wire \onchip_memory2_0_s1_writedata[8]~input_o ;
wire \onchip_memory2_0_s1_byteenable[1]~input_o ;
wire \onchip_memory2_0_s2_writedata[8]~input_o ;
wire \onchip_memory2_0_s2_byteenable[1]~input_o ;
wire \onchip_memory2_0_s1_writedata[9]~input_o ;
wire \onchip_memory2_0_s2_writedata[9]~input_o ;
wire \onchip_memory2_0_s1_writedata[10]~input_o ;
wire \onchip_memory2_0_s2_writedata[10]~input_o ;
wire \onchip_memory2_0_s1_writedata[11]~input_o ;
wire \onchip_memory2_0_s2_writedata[11]~input_o ;
wire \onchip_memory2_0_s1_writedata[12]~input_o ;
wire \onchip_memory2_0_s2_writedata[12]~input_o ;
wire \onchip_memory2_0_s1_writedata[13]~input_o ;
wire \onchip_memory2_0_s2_writedata[13]~input_o ;
wire \onchip_memory2_0_s1_writedata[14]~input_o ;
wire \onchip_memory2_0_s2_writedata[14]~input_o ;
wire \onchip_memory2_0_s1_writedata[15]~input_o ;
wire \onchip_memory2_0_s2_writedata[15]~input_o ;
wire \onchip_memory2_0_s1_writedata[16]~input_o ;
wire \onchip_memory2_0_s1_byteenable[2]~input_o ;
wire \onchip_memory2_0_s2_writedata[16]~input_o ;
wire \onchip_memory2_0_s2_byteenable[2]~input_o ;
wire \onchip_memory2_0_s1_writedata[17]~input_o ;
wire \onchip_memory2_0_s2_writedata[17]~input_o ;
wire \onchip_memory2_0_s1_writedata[18]~input_o ;
wire \onchip_memory2_0_s2_writedata[18]~input_o ;
wire \onchip_memory2_0_s1_writedata[19]~input_o ;
wire \onchip_memory2_0_s2_writedata[19]~input_o ;
wire \onchip_memory2_0_s1_writedata[20]~input_o ;
wire \onchip_memory2_0_s2_writedata[20]~input_o ;
wire \onchip_memory2_0_s1_writedata[21]~input_o ;
wire \onchip_memory2_0_s2_writedata[21]~input_o ;
wire \onchip_memory2_0_s1_writedata[22]~input_o ;
wire \onchip_memory2_0_s2_writedata[22]~input_o ;
wire \onchip_memory2_0_s1_writedata[23]~input_o ;
wire \onchip_memory2_0_s2_writedata[23]~input_o ;
wire \onchip_memory2_0_s1_writedata[24]~input_o ;
wire \onchip_memory2_0_s1_byteenable[3]~input_o ;
wire \onchip_memory2_0_s2_writedata[24]~input_o ;
wire \onchip_memory2_0_s2_byteenable[3]~input_o ;
wire \onchip_memory2_0_s1_writedata[25]~input_o ;
wire \onchip_memory2_0_s2_writedata[25]~input_o ;
wire \onchip_memory2_0_s1_writedata[26]~input_o ;
wire \onchip_memory2_0_s2_writedata[26]~input_o ;
wire \onchip_memory2_0_s1_writedata[27]~input_o ;
wire \onchip_memory2_0_s2_writedata[27]~input_o ;
wire \onchip_memory2_0_s1_writedata[28]~input_o ;
wire \onchip_memory2_0_s2_writedata[28]~input_o ;
wire \onchip_memory2_0_s1_writedata[29]~input_o ;
wire \onchip_memory2_0_s2_writedata[29]~input_o ;
wire \onchip_memory2_0_s1_writedata[30]~input_o ;
wire \onchip_memory2_0_s2_writedata[30]~input_o ;
wire \onchip_memory2_0_s1_writedata[31]~input_o ;
wire \onchip_memory2_0_s2_writedata[31]~input_o ;
wire \onchip_memory2_0_s1_writedata[32]~input_o ;
wire \onchip_memory2_0_s1_byteenable[4]~input_o ;
wire \onchip_memory2_0_s2_writedata[32]~input_o ;
wire \onchip_memory2_0_s2_byteenable[4]~input_o ;
wire \onchip_memory2_0_s1_writedata[33]~input_o ;
wire \onchip_memory2_0_s2_writedata[33]~input_o ;
wire \onchip_memory2_0_s1_writedata[34]~input_o ;
wire \onchip_memory2_0_s2_writedata[34]~input_o ;
wire \onchip_memory2_0_s1_writedata[35]~input_o ;
wire \onchip_memory2_0_s2_writedata[35]~input_o ;
wire \onchip_memory2_0_s1_writedata[36]~input_o ;
wire \onchip_memory2_0_s2_writedata[36]~input_o ;
wire \onchip_memory2_0_s1_writedata[37]~input_o ;
wire \onchip_memory2_0_s2_writedata[37]~input_o ;
wire \onchip_memory2_0_s1_writedata[38]~input_o ;
wire \onchip_memory2_0_s2_writedata[38]~input_o ;
wire \onchip_memory2_0_s1_writedata[39]~input_o ;
wire \onchip_memory2_0_s2_writedata[39]~input_o ;
wire \onchip_memory2_0_s1_writedata[40]~input_o ;
wire \onchip_memory2_0_s1_byteenable[5]~input_o ;
wire \onchip_memory2_0_s2_writedata[40]~input_o ;
wire \onchip_memory2_0_s2_byteenable[5]~input_o ;
wire \onchip_memory2_0_s1_writedata[41]~input_o ;
wire \onchip_memory2_0_s2_writedata[41]~input_o ;
wire \onchip_memory2_0_s1_writedata[42]~input_o ;
wire \onchip_memory2_0_s2_writedata[42]~input_o ;
wire \onchip_memory2_0_s1_writedata[43]~input_o ;
wire \onchip_memory2_0_s2_writedata[43]~input_o ;
wire \onchip_memory2_0_s1_writedata[44]~input_o ;
wire \onchip_memory2_0_s2_writedata[44]~input_o ;
wire \onchip_memory2_0_s1_writedata[45]~input_o ;
wire \onchip_memory2_0_s2_writedata[45]~input_o ;
wire \onchip_memory2_0_s1_writedata[46]~input_o ;
wire \onchip_memory2_0_s2_writedata[46]~input_o ;
wire \onchip_memory2_0_s1_writedata[47]~input_o ;
wire \onchip_memory2_0_s2_writedata[47]~input_o ;
wire \onchip_memory2_0_s1_writedata[48]~input_o ;
wire \onchip_memory2_0_s1_byteenable[6]~input_o ;
wire \onchip_memory2_0_s2_writedata[48]~input_o ;
wire \onchip_memory2_0_s2_byteenable[6]~input_o ;
wire \onchip_memory2_0_s1_writedata[49]~input_o ;
wire \onchip_memory2_0_s2_writedata[49]~input_o ;
wire \onchip_memory2_0_s1_writedata[50]~input_o ;
wire \onchip_memory2_0_s2_writedata[50]~input_o ;
wire \onchip_memory2_0_s1_writedata[51]~input_o ;
wire \onchip_memory2_0_s2_writedata[51]~input_o ;
wire \onchip_memory2_0_s1_writedata[52]~input_o ;
wire \onchip_memory2_0_s2_writedata[52]~input_o ;
wire \onchip_memory2_0_s1_writedata[53]~input_o ;
wire \onchip_memory2_0_s2_writedata[53]~input_o ;
wire \onchip_memory2_0_s1_writedata[54]~input_o ;
wire \onchip_memory2_0_s2_writedata[54]~input_o ;
wire \onchip_memory2_0_s1_writedata[55]~input_o ;
wire \onchip_memory2_0_s2_writedata[55]~input_o ;
wire \onchip_memory2_0_s1_writedata[56]~input_o ;
wire \onchip_memory2_0_s1_byteenable[7]~input_o ;
wire \onchip_memory2_0_s2_writedata[56]~input_o ;
wire \onchip_memory2_0_s2_byteenable[7]~input_o ;
wire \onchip_memory2_0_s1_writedata[57]~input_o ;
wire \onchip_memory2_0_s2_writedata[57]~input_o ;
wire \onchip_memory2_0_s1_writedata[58]~input_o ;
wire \onchip_memory2_0_s2_writedata[58]~input_o ;
wire \onchip_memory2_0_s1_writedata[59]~input_o ;
wire \onchip_memory2_0_s2_writedata[59]~input_o ;
wire \onchip_memory2_0_s1_writedata[60]~input_o ;
wire \onchip_memory2_0_s2_writedata[60]~input_o ;
wire \onchip_memory2_0_s1_writedata[61]~input_o ;
wire \onchip_memory2_0_s2_writedata[61]~input_o ;
wire \onchip_memory2_0_s1_writedata[62]~input_o ;
wire \onchip_memory2_0_s2_writedata[62]~input_o ;
wire \onchip_memory2_0_s1_writedata[63]~input_o ;
wire \onchip_memory2_0_s2_writedata[63]~input_o ;
wire \reset_reset_n~input_o ;


qtestpd_altera_reset_controller rst_controller(
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.clk_clk(\clk_clk~input_o ),
	.reset_reset_n(\reset_reset_n~input_o ));

qtestpd_qtestpd_onchip_memory2_0 onchip_memory2_0(
	.result_node_0(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[0]~0_combout ),
	.result_node_1(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[1]~1_combout ),
	.result_node_2(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[2]~2_combout ),
	.result_node_3(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[3]~3_combout ),
	.result_node_4(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[4]~4_combout ),
	.result_node_5(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[5]~5_combout ),
	.result_node_6(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[6]~6_combout ),
	.result_node_7(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[7]~7_combout ),
	.result_node_8(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[8]~8_combout ),
	.result_node_9(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[9]~9_combout ),
	.result_node_10(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[10]~10_combout ),
	.result_node_11(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[11]~11_combout ),
	.result_node_12(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[12]~12_combout ),
	.result_node_13(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[13]~13_combout ),
	.result_node_14(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[14]~14_combout ),
	.result_node_15(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[15]~15_combout ),
	.result_node_16(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[16]~16_combout ),
	.result_node_17(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[17]~17_combout ),
	.result_node_18(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[18]~18_combout ),
	.result_node_19(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[19]~19_combout ),
	.result_node_20(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[20]~20_combout ),
	.result_node_21(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[21]~21_combout ),
	.result_node_22(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[22]~22_combout ),
	.result_node_23(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[23]~23_combout ),
	.result_node_24(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[24]~24_combout ),
	.result_node_25(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[25]~25_combout ),
	.result_node_26(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[26]~26_combout ),
	.result_node_27(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[27]~27_combout ),
	.result_node_28(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[28]~28_combout ),
	.result_node_29(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[29]~29_combout ),
	.result_node_30(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[30]~30_combout ),
	.result_node_31(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[31]~31_combout ),
	.result_node_32(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[32]~32_combout ),
	.result_node_33(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[33]~33_combout ),
	.result_node_34(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[34]~34_combout ),
	.result_node_35(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[35]~35_combout ),
	.result_node_36(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[36]~36_combout ),
	.result_node_37(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[37]~37_combout ),
	.result_node_38(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[38]~38_combout ),
	.result_node_39(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[39]~39_combout ),
	.result_node_40(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[40]~40_combout ),
	.result_node_41(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[41]~41_combout ),
	.result_node_42(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[42]~42_combout ),
	.result_node_43(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[43]~43_combout ),
	.result_node_44(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[44]~44_combout ),
	.result_node_45(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[45]~45_combout ),
	.result_node_46(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[46]~46_combout ),
	.result_node_47(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[47]~47_combout ),
	.result_node_48(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[48]~48_combout ),
	.result_node_49(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[49]~49_combout ),
	.result_node_50(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[50]~50_combout ),
	.result_node_51(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[51]~51_combout ),
	.result_node_52(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[52]~52_combout ),
	.result_node_53(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[53]~53_combout ),
	.result_node_54(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[54]~54_combout ),
	.result_node_55(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[55]~55_combout ),
	.result_node_56(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[56]~56_combout ),
	.result_node_57(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[57]~57_combout ),
	.result_node_58(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[58]~58_combout ),
	.result_node_59(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[59]~59_combout ),
	.result_node_60(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[60]~60_combout ),
	.result_node_61(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[61]~61_combout ),
	.result_node_62(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[62]~62_combout ),
	.result_node_63(\onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[63]~63_combout ),
	.result_node_01(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[0]~0_combout ),
	.result_node_110(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[1]~1_combout ),
	.result_node_210(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[2]~2_combout ),
	.result_node_310(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[3]~3_combout ),
	.result_node_410(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[4]~4_combout ),
	.result_node_510(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[5]~5_combout ),
	.result_node_64(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[6]~6_combout ),
	.result_node_71(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[7]~7_combout ),
	.result_node_81(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[8]~8_combout ),
	.result_node_91(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[9]~9_combout ),
	.result_node_101(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[10]~10_combout ),
	.result_node_111(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[11]~11_combout ),
	.result_node_121(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[12]~12_combout ),
	.result_node_131(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[13]~13_combout ),
	.result_node_141(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[14]~14_combout ),
	.result_node_151(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[15]~15_combout ),
	.result_node_161(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[16]~16_combout ),
	.result_node_171(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[17]~17_combout ),
	.result_node_181(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[18]~18_combout ),
	.result_node_191(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[19]~19_combout ),
	.result_node_201(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[20]~20_combout ),
	.result_node_211(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[21]~21_combout ),
	.result_node_221(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[22]~22_combout ),
	.result_node_231(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[23]~23_combout ),
	.result_node_241(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[24]~24_combout ),
	.result_node_251(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[25]~25_combout ),
	.result_node_261(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[26]~26_combout ),
	.result_node_271(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[27]~27_combout ),
	.result_node_281(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[28]~28_combout ),
	.result_node_291(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[29]~29_combout ),
	.result_node_301(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[30]~30_combout ),
	.result_node_311(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[31]~31_combout ),
	.result_node_321(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[32]~32_combout ),
	.result_node_331(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[33]~33_combout ),
	.result_node_341(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[34]~34_combout ),
	.result_node_351(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[35]~35_combout ),
	.result_node_361(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[36]~36_combout ),
	.result_node_371(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[37]~37_combout ),
	.result_node_381(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[38]~38_combout ),
	.result_node_391(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[39]~39_combout ),
	.result_node_401(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[40]~40_combout ),
	.result_node_411(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[41]~41_combout ),
	.result_node_421(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[42]~42_combout ),
	.result_node_431(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[43]~43_combout ),
	.result_node_441(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[44]~44_combout ),
	.result_node_451(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[45]~45_combout ),
	.result_node_461(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[46]~46_combout ),
	.result_node_471(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[47]~47_combout ),
	.result_node_481(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[48]~48_combout ),
	.result_node_491(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[49]~49_combout ),
	.result_node_501(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[50]~50_combout ),
	.result_node_511(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[51]~51_combout ),
	.result_node_521(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[52]~52_combout ),
	.result_node_531(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[53]~53_combout ),
	.result_node_541(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[54]~54_combout ),
	.result_node_551(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[55]~55_combout ),
	.result_node_561(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[56]~56_combout ),
	.result_node_571(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[57]~57_combout ),
	.result_node_581(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[58]~58_combout ),
	.result_node_591(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[59]~59_combout ),
	.result_node_601(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[60]~60_combout ),
	.result_node_611(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[61]~61_combout ),
	.result_node_621(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[62]~62_combout ),
	.result_node_631(\onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[63]~63_combout ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.onchip_memory2_0_s1_address_13(\onchip_memory2_0_s1_address[13]~input_o ),
	.onchip_memory2_0_s1_chipselect(\onchip_memory2_0_s1_chipselect~input_o ),
	.onchip_memory2_0_s1_write(\onchip_memory2_0_s1_write~input_o ),
	.onchip_memory2_0_s2_address_13(\onchip_memory2_0_s2_address[13]~input_o ),
	.onchip_memory2_0_s2_chipselect(\onchip_memory2_0_s2_chipselect~input_o ),
	.onchip_memory2_0_s2_write(\onchip_memory2_0_s2_write~input_o ),
	.clk_clk(\clk_clk~input_o ),
	.onchip_memory2_0_s1_clken(\onchip_memory2_0_s1_clken~input_o ),
	.onchip_memory2_0_s2_clken(\onchip_memory2_0_s2_clken~input_o ),
	.onchip_memory2_0_s1_writedata_0(\onchip_memory2_0_s1_writedata[0]~input_o ),
	.onchip_memory2_0_s1_address_0(\onchip_memory2_0_s1_address[0]~input_o ),
	.onchip_memory2_0_s1_address_1(\onchip_memory2_0_s1_address[1]~input_o ),
	.onchip_memory2_0_s1_address_2(\onchip_memory2_0_s1_address[2]~input_o ),
	.onchip_memory2_0_s1_address_3(\onchip_memory2_0_s1_address[3]~input_o ),
	.onchip_memory2_0_s1_address_4(\onchip_memory2_0_s1_address[4]~input_o ),
	.onchip_memory2_0_s1_address_5(\onchip_memory2_0_s1_address[5]~input_o ),
	.onchip_memory2_0_s1_address_6(\onchip_memory2_0_s1_address[6]~input_o ),
	.onchip_memory2_0_s1_address_7(\onchip_memory2_0_s1_address[7]~input_o ),
	.onchip_memory2_0_s1_address_8(\onchip_memory2_0_s1_address[8]~input_o ),
	.onchip_memory2_0_s1_address_9(\onchip_memory2_0_s1_address[9]~input_o ),
	.onchip_memory2_0_s1_address_10(\onchip_memory2_0_s1_address[10]~input_o ),
	.onchip_memory2_0_s1_address_11(\onchip_memory2_0_s1_address[11]~input_o ),
	.onchip_memory2_0_s1_address_12(\onchip_memory2_0_s1_address[12]~input_o ),
	.onchip_memory2_0_s1_byteenable_0(\onchip_memory2_0_s1_byteenable[0]~input_o ),
	.onchip_memory2_0_s2_writedata_0(\onchip_memory2_0_s2_writedata[0]~input_o ),
	.onchip_memory2_0_s2_address_0(\onchip_memory2_0_s2_address[0]~input_o ),
	.onchip_memory2_0_s2_address_1(\onchip_memory2_0_s2_address[1]~input_o ),
	.onchip_memory2_0_s2_address_2(\onchip_memory2_0_s2_address[2]~input_o ),
	.onchip_memory2_0_s2_address_3(\onchip_memory2_0_s2_address[3]~input_o ),
	.onchip_memory2_0_s2_address_4(\onchip_memory2_0_s2_address[4]~input_o ),
	.onchip_memory2_0_s2_address_5(\onchip_memory2_0_s2_address[5]~input_o ),
	.onchip_memory2_0_s2_address_6(\onchip_memory2_0_s2_address[6]~input_o ),
	.onchip_memory2_0_s2_address_7(\onchip_memory2_0_s2_address[7]~input_o ),
	.onchip_memory2_0_s2_address_8(\onchip_memory2_0_s2_address[8]~input_o ),
	.onchip_memory2_0_s2_address_9(\onchip_memory2_0_s2_address[9]~input_o ),
	.onchip_memory2_0_s2_address_10(\onchip_memory2_0_s2_address[10]~input_o ),
	.onchip_memory2_0_s2_address_11(\onchip_memory2_0_s2_address[11]~input_o ),
	.onchip_memory2_0_s2_address_12(\onchip_memory2_0_s2_address[12]~input_o ),
	.onchip_memory2_0_s2_byteenable_0(\onchip_memory2_0_s2_byteenable[0]~input_o ),
	.onchip_memory2_0_s1_writedata_1(\onchip_memory2_0_s1_writedata[1]~input_o ),
	.onchip_memory2_0_s2_writedata_1(\onchip_memory2_0_s2_writedata[1]~input_o ),
	.onchip_memory2_0_s1_writedata_2(\onchip_memory2_0_s1_writedata[2]~input_o ),
	.onchip_memory2_0_s2_writedata_2(\onchip_memory2_0_s2_writedata[2]~input_o ),
	.onchip_memory2_0_s1_writedata_3(\onchip_memory2_0_s1_writedata[3]~input_o ),
	.onchip_memory2_0_s2_writedata_3(\onchip_memory2_0_s2_writedata[3]~input_o ),
	.onchip_memory2_0_s1_writedata_4(\onchip_memory2_0_s1_writedata[4]~input_o ),
	.onchip_memory2_0_s2_writedata_4(\onchip_memory2_0_s2_writedata[4]~input_o ),
	.onchip_memory2_0_s1_writedata_5(\onchip_memory2_0_s1_writedata[5]~input_o ),
	.onchip_memory2_0_s2_writedata_5(\onchip_memory2_0_s2_writedata[5]~input_o ),
	.onchip_memory2_0_s1_writedata_6(\onchip_memory2_0_s1_writedata[6]~input_o ),
	.onchip_memory2_0_s2_writedata_6(\onchip_memory2_0_s2_writedata[6]~input_o ),
	.onchip_memory2_0_s1_writedata_7(\onchip_memory2_0_s1_writedata[7]~input_o ),
	.onchip_memory2_0_s2_writedata_7(\onchip_memory2_0_s2_writedata[7]~input_o ),
	.onchip_memory2_0_s1_writedata_8(\onchip_memory2_0_s1_writedata[8]~input_o ),
	.onchip_memory2_0_s1_byteenable_1(\onchip_memory2_0_s1_byteenable[1]~input_o ),
	.onchip_memory2_0_s2_writedata_8(\onchip_memory2_0_s2_writedata[8]~input_o ),
	.onchip_memory2_0_s2_byteenable_1(\onchip_memory2_0_s2_byteenable[1]~input_o ),
	.onchip_memory2_0_s1_writedata_9(\onchip_memory2_0_s1_writedata[9]~input_o ),
	.onchip_memory2_0_s2_writedata_9(\onchip_memory2_0_s2_writedata[9]~input_o ),
	.onchip_memory2_0_s1_writedata_10(\onchip_memory2_0_s1_writedata[10]~input_o ),
	.onchip_memory2_0_s2_writedata_10(\onchip_memory2_0_s2_writedata[10]~input_o ),
	.onchip_memory2_0_s1_writedata_11(\onchip_memory2_0_s1_writedata[11]~input_o ),
	.onchip_memory2_0_s2_writedata_11(\onchip_memory2_0_s2_writedata[11]~input_o ),
	.onchip_memory2_0_s1_writedata_12(\onchip_memory2_0_s1_writedata[12]~input_o ),
	.onchip_memory2_0_s2_writedata_12(\onchip_memory2_0_s2_writedata[12]~input_o ),
	.onchip_memory2_0_s1_writedata_13(\onchip_memory2_0_s1_writedata[13]~input_o ),
	.onchip_memory2_0_s2_writedata_13(\onchip_memory2_0_s2_writedata[13]~input_o ),
	.onchip_memory2_0_s1_writedata_14(\onchip_memory2_0_s1_writedata[14]~input_o ),
	.onchip_memory2_0_s2_writedata_14(\onchip_memory2_0_s2_writedata[14]~input_o ),
	.onchip_memory2_0_s1_writedata_15(\onchip_memory2_0_s1_writedata[15]~input_o ),
	.onchip_memory2_0_s2_writedata_15(\onchip_memory2_0_s2_writedata[15]~input_o ),
	.onchip_memory2_0_s1_writedata_16(\onchip_memory2_0_s1_writedata[16]~input_o ),
	.onchip_memory2_0_s1_byteenable_2(\onchip_memory2_0_s1_byteenable[2]~input_o ),
	.onchip_memory2_0_s2_writedata_16(\onchip_memory2_0_s2_writedata[16]~input_o ),
	.onchip_memory2_0_s2_byteenable_2(\onchip_memory2_0_s2_byteenable[2]~input_o ),
	.onchip_memory2_0_s1_writedata_17(\onchip_memory2_0_s1_writedata[17]~input_o ),
	.onchip_memory2_0_s2_writedata_17(\onchip_memory2_0_s2_writedata[17]~input_o ),
	.onchip_memory2_0_s1_writedata_18(\onchip_memory2_0_s1_writedata[18]~input_o ),
	.onchip_memory2_0_s2_writedata_18(\onchip_memory2_0_s2_writedata[18]~input_o ),
	.onchip_memory2_0_s1_writedata_19(\onchip_memory2_0_s1_writedata[19]~input_o ),
	.onchip_memory2_0_s2_writedata_19(\onchip_memory2_0_s2_writedata[19]~input_o ),
	.onchip_memory2_0_s1_writedata_20(\onchip_memory2_0_s1_writedata[20]~input_o ),
	.onchip_memory2_0_s2_writedata_20(\onchip_memory2_0_s2_writedata[20]~input_o ),
	.onchip_memory2_0_s1_writedata_21(\onchip_memory2_0_s1_writedata[21]~input_o ),
	.onchip_memory2_0_s2_writedata_21(\onchip_memory2_0_s2_writedata[21]~input_o ),
	.onchip_memory2_0_s1_writedata_22(\onchip_memory2_0_s1_writedata[22]~input_o ),
	.onchip_memory2_0_s2_writedata_22(\onchip_memory2_0_s2_writedata[22]~input_o ),
	.onchip_memory2_0_s1_writedata_23(\onchip_memory2_0_s1_writedata[23]~input_o ),
	.onchip_memory2_0_s2_writedata_23(\onchip_memory2_0_s2_writedata[23]~input_o ),
	.onchip_memory2_0_s1_writedata_24(\onchip_memory2_0_s1_writedata[24]~input_o ),
	.onchip_memory2_0_s1_byteenable_3(\onchip_memory2_0_s1_byteenable[3]~input_o ),
	.onchip_memory2_0_s2_writedata_24(\onchip_memory2_0_s2_writedata[24]~input_o ),
	.onchip_memory2_0_s2_byteenable_3(\onchip_memory2_0_s2_byteenable[3]~input_o ),
	.onchip_memory2_0_s1_writedata_25(\onchip_memory2_0_s1_writedata[25]~input_o ),
	.onchip_memory2_0_s2_writedata_25(\onchip_memory2_0_s2_writedata[25]~input_o ),
	.onchip_memory2_0_s1_writedata_26(\onchip_memory2_0_s1_writedata[26]~input_o ),
	.onchip_memory2_0_s2_writedata_26(\onchip_memory2_0_s2_writedata[26]~input_o ),
	.onchip_memory2_0_s1_writedata_27(\onchip_memory2_0_s1_writedata[27]~input_o ),
	.onchip_memory2_0_s2_writedata_27(\onchip_memory2_0_s2_writedata[27]~input_o ),
	.onchip_memory2_0_s1_writedata_28(\onchip_memory2_0_s1_writedata[28]~input_o ),
	.onchip_memory2_0_s2_writedata_28(\onchip_memory2_0_s2_writedata[28]~input_o ),
	.onchip_memory2_0_s1_writedata_29(\onchip_memory2_0_s1_writedata[29]~input_o ),
	.onchip_memory2_0_s2_writedata_29(\onchip_memory2_0_s2_writedata[29]~input_o ),
	.onchip_memory2_0_s1_writedata_30(\onchip_memory2_0_s1_writedata[30]~input_o ),
	.onchip_memory2_0_s2_writedata_30(\onchip_memory2_0_s2_writedata[30]~input_o ),
	.onchip_memory2_0_s1_writedata_31(\onchip_memory2_0_s1_writedata[31]~input_o ),
	.onchip_memory2_0_s2_writedata_31(\onchip_memory2_0_s2_writedata[31]~input_o ),
	.onchip_memory2_0_s1_writedata_32(\onchip_memory2_0_s1_writedata[32]~input_o ),
	.onchip_memory2_0_s1_byteenable_4(\onchip_memory2_0_s1_byteenable[4]~input_o ),
	.onchip_memory2_0_s2_writedata_32(\onchip_memory2_0_s2_writedata[32]~input_o ),
	.onchip_memory2_0_s2_byteenable_4(\onchip_memory2_0_s2_byteenable[4]~input_o ),
	.onchip_memory2_0_s1_writedata_33(\onchip_memory2_0_s1_writedata[33]~input_o ),
	.onchip_memory2_0_s2_writedata_33(\onchip_memory2_0_s2_writedata[33]~input_o ),
	.onchip_memory2_0_s1_writedata_34(\onchip_memory2_0_s1_writedata[34]~input_o ),
	.onchip_memory2_0_s2_writedata_34(\onchip_memory2_0_s2_writedata[34]~input_o ),
	.onchip_memory2_0_s1_writedata_35(\onchip_memory2_0_s1_writedata[35]~input_o ),
	.onchip_memory2_0_s2_writedata_35(\onchip_memory2_0_s2_writedata[35]~input_o ),
	.onchip_memory2_0_s1_writedata_36(\onchip_memory2_0_s1_writedata[36]~input_o ),
	.onchip_memory2_0_s2_writedata_36(\onchip_memory2_0_s2_writedata[36]~input_o ),
	.onchip_memory2_0_s1_writedata_37(\onchip_memory2_0_s1_writedata[37]~input_o ),
	.onchip_memory2_0_s2_writedata_37(\onchip_memory2_0_s2_writedata[37]~input_o ),
	.onchip_memory2_0_s1_writedata_38(\onchip_memory2_0_s1_writedata[38]~input_o ),
	.onchip_memory2_0_s2_writedata_38(\onchip_memory2_0_s2_writedata[38]~input_o ),
	.onchip_memory2_0_s1_writedata_39(\onchip_memory2_0_s1_writedata[39]~input_o ),
	.onchip_memory2_0_s2_writedata_39(\onchip_memory2_0_s2_writedata[39]~input_o ),
	.onchip_memory2_0_s1_writedata_40(\onchip_memory2_0_s1_writedata[40]~input_o ),
	.onchip_memory2_0_s1_byteenable_5(\onchip_memory2_0_s1_byteenable[5]~input_o ),
	.onchip_memory2_0_s2_writedata_40(\onchip_memory2_0_s2_writedata[40]~input_o ),
	.onchip_memory2_0_s2_byteenable_5(\onchip_memory2_0_s2_byteenable[5]~input_o ),
	.onchip_memory2_0_s1_writedata_41(\onchip_memory2_0_s1_writedata[41]~input_o ),
	.onchip_memory2_0_s2_writedata_41(\onchip_memory2_0_s2_writedata[41]~input_o ),
	.onchip_memory2_0_s1_writedata_42(\onchip_memory2_0_s1_writedata[42]~input_o ),
	.onchip_memory2_0_s2_writedata_42(\onchip_memory2_0_s2_writedata[42]~input_o ),
	.onchip_memory2_0_s1_writedata_43(\onchip_memory2_0_s1_writedata[43]~input_o ),
	.onchip_memory2_0_s2_writedata_43(\onchip_memory2_0_s2_writedata[43]~input_o ),
	.onchip_memory2_0_s1_writedata_44(\onchip_memory2_0_s1_writedata[44]~input_o ),
	.onchip_memory2_0_s2_writedata_44(\onchip_memory2_0_s2_writedata[44]~input_o ),
	.onchip_memory2_0_s1_writedata_45(\onchip_memory2_0_s1_writedata[45]~input_o ),
	.onchip_memory2_0_s2_writedata_45(\onchip_memory2_0_s2_writedata[45]~input_o ),
	.onchip_memory2_0_s1_writedata_46(\onchip_memory2_0_s1_writedata[46]~input_o ),
	.onchip_memory2_0_s2_writedata_46(\onchip_memory2_0_s2_writedata[46]~input_o ),
	.onchip_memory2_0_s1_writedata_47(\onchip_memory2_0_s1_writedata[47]~input_o ),
	.onchip_memory2_0_s2_writedata_47(\onchip_memory2_0_s2_writedata[47]~input_o ),
	.onchip_memory2_0_s1_writedata_48(\onchip_memory2_0_s1_writedata[48]~input_o ),
	.onchip_memory2_0_s1_byteenable_6(\onchip_memory2_0_s1_byteenable[6]~input_o ),
	.onchip_memory2_0_s2_writedata_48(\onchip_memory2_0_s2_writedata[48]~input_o ),
	.onchip_memory2_0_s2_byteenable_6(\onchip_memory2_0_s2_byteenable[6]~input_o ),
	.onchip_memory2_0_s1_writedata_49(\onchip_memory2_0_s1_writedata[49]~input_o ),
	.onchip_memory2_0_s2_writedata_49(\onchip_memory2_0_s2_writedata[49]~input_o ),
	.onchip_memory2_0_s1_writedata_50(\onchip_memory2_0_s1_writedata[50]~input_o ),
	.onchip_memory2_0_s2_writedata_50(\onchip_memory2_0_s2_writedata[50]~input_o ),
	.onchip_memory2_0_s1_writedata_51(\onchip_memory2_0_s1_writedata[51]~input_o ),
	.onchip_memory2_0_s2_writedata_51(\onchip_memory2_0_s2_writedata[51]~input_o ),
	.onchip_memory2_0_s1_writedata_52(\onchip_memory2_0_s1_writedata[52]~input_o ),
	.onchip_memory2_0_s2_writedata_52(\onchip_memory2_0_s2_writedata[52]~input_o ),
	.onchip_memory2_0_s1_writedata_53(\onchip_memory2_0_s1_writedata[53]~input_o ),
	.onchip_memory2_0_s2_writedata_53(\onchip_memory2_0_s2_writedata[53]~input_o ),
	.onchip_memory2_0_s1_writedata_54(\onchip_memory2_0_s1_writedata[54]~input_o ),
	.onchip_memory2_0_s2_writedata_54(\onchip_memory2_0_s2_writedata[54]~input_o ),
	.onchip_memory2_0_s1_writedata_55(\onchip_memory2_0_s1_writedata[55]~input_o ),
	.onchip_memory2_0_s2_writedata_55(\onchip_memory2_0_s2_writedata[55]~input_o ),
	.onchip_memory2_0_s1_writedata_56(\onchip_memory2_0_s1_writedata[56]~input_o ),
	.onchip_memory2_0_s1_byteenable_7(\onchip_memory2_0_s1_byteenable[7]~input_o ),
	.onchip_memory2_0_s2_writedata_56(\onchip_memory2_0_s2_writedata[56]~input_o ),
	.onchip_memory2_0_s2_byteenable_7(\onchip_memory2_0_s2_byteenable[7]~input_o ),
	.onchip_memory2_0_s1_writedata_57(\onchip_memory2_0_s1_writedata[57]~input_o ),
	.onchip_memory2_0_s2_writedata_57(\onchip_memory2_0_s2_writedata[57]~input_o ),
	.onchip_memory2_0_s1_writedata_58(\onchip_memory2_0_s1_writedata[58]~input_o ),
	.onchip_memory2_0_s2_writedata_58(\onchip_memory2_0_s2_writedata[58]~input_o ),
	.onchip_memory2_0_s1_writedata_59(\onchip_memory2_0_s1_writedata[59]~input_o ),
	.onchip_memory2_0_s2_writedata_59(\onchip_memory2_0_s2_writedata[59]~input_o ),
	.onchip_memory2_0_s1_writedata_60(\onchip_memory2_0_s1_writedata[60]~input_o ),
	.onchip_memory2_0_s2_writedata_60(\onchip_memory2_0_s2_writedata[60]~input_o ),
	.onchip_memory2_0_s1_writedata_61(\onchip_memory2_0_s1_writedata[61]~input_o ),
	.onchip_memory2_0_s2_writedata_61(\onchip_memory2_0_s2_writedata[61]~input_o ),
	.onchip_memory2_0_s1_writedata_62(\onchip_memory2_0_s1_writedata[62]~input_o ),
	.onchip_memory2_0_s2_writedata_62(\onchip_memory2_0_s2_writedata[62]~input_o ),
	.onchip_memory2_0_s1_writedata_63(\onchip_memory2_0_s1_writedata[63]~input_o ),
	.onchip_memory2_0_s2_writedata_63(\onchip_memory2_0_s2_writedata[63]~input_o ));

assign \onchip_memory2_0_s1_address[13]~input_o  = onchip_memory2_0_s1_address[13];

assign \onchip_memory2_0_s1_chipselect~input_o  = onchip_memory2_0_s1_chipselect;

assign \onchip_memory2_0_s1_write~input_o  = onchip_memory2_0_s1_write;

assign \onchip_memory2_0_s2_address[13]~input_o  = onchip_memory2_0_s2_address[13];

assign \onchip_memory2_0_s2_chipselect~input_o  = onchip_memory2_0_s2_chipselect;

assign \onchip_memory2_0_s2_write~input_o  = onchip_memory2_0_s2_write;

assign \clk_clk~input_o  = clk_clk;

assign \onchip_memory2_0_s1_clken~input_o  = onchip_memory2_0_s1_clken;

assign \onchip_memory2_0_s2_clken~input_o  = onchip_memory2_0_s2_clken;

assign \onchip_memory2_0_s1_writedata[0]~input_o  = onchip_memory2_0_s1_writedata[0];

assign \onchip_memory2_0_s1_address[0]~input_o  = onchip_memory2_0_s1_address[0];

assign \onchip_memory2_0_s1_address[1]~input_o  = onchip_memory2_0_s1_address[1];

assign \onchip_memory2_0_s1_address[2]~input_o  = onchip_memory2_0_s1_address[2];

assign \onchip_memory2_0_s1_address[3]~input_o  = onchip_memory2_0_s1_address[3];

assign \onchip_memory2_0_s1_address[4]~input_o  = onchip_memory2_0_s1_address[4];

assign \onchip_memory2_0_s1_address[5]~input_o  = onchip_memory2_0_s1_address[5];

assign \onchip_memory2_0_s1_address[6]~input_o  = onchip_memory2_0_s1_address[6];

assign \onchip_memory2_0_s1_address[7]~input_o  = onchip_memory2_0_s1_address[7];

assign \onchip_memory2_0_s1_address[8]~input_o  = onchip_memory2_0_s1_address[8];

assign \onchip_memory2_0_s1_address[9]~input_o  = onchip_memory2_0_s1_address[9];

assign \onchip_memory2_0_s1_address[10]~input_o  = onchip_memory2_0_s1_address[10];

assign \onchip_memory2_0_s1_address[11]~input_o  = onchip_memory2_0_s1_address[11];

assign \onchip_memory2_0_s1_address[12]~input_o  = onchip_memory2_0_s1_address[12];

assign \onchip_memory2_0_s1_byteenable[0]~input_o  = onchip_memory2_0_s1_byteenable[0];

assign \onchip_memory2_0_s2_writedata[0]~input_o  = onchip_memory2_0_s2_writedata[0];

assign \onchip_memory2_0_s2_address[0]~input_o  = onchip_memory2_0_s2_address[0];

assign \onchip_memory2_0_s2_address[1]~input_o  = onchip_memory2_0_s2_address[1];

assign \onchip_memory2_0_s2_address[2]~input_o  = onchip_memory2_0_s2_address[2];

assign \onchip_memory2_0_s2_address[3]~input_o  = onchip_memory2_0_s2_address[3];

assign \onchip_memory2_0_s2_address[4]~input_o  = onchip_memory2_0_s2_address[4];

assign \onchip_memory2_0_s2_address[5]~input_o  = onchip_memory2_0_s2_address[5];

assign \onchip_memory2_0_s2_address[6]~input_o  = onchip_memory2_0_s2_address[6];

assign \onchip_memory2_0_s2_address[7]~input_o  = onchip_memory2_0_s2_address[7];

assign \onchip_memory2_0_s2_address[8]~input_o  = onchip_memory2_0_s2_address[8];

assign \onchip_memory2_0_s2_address[9]~input_o  = onchip_memory2_0_s2_address[9];

assign \onchip_memory2_0_s2_address[10]~input_o  = onchip_memory2_0_s2_address[10];

assign \onchip_memory2_0_s2_address[11]~input_o  = onchip_memory2_0_s2_address[11];

assign \onchip_memory2_0_s2_address[12]~input_o  = onchip_memory2_0_s2_address[12];

assign \onchip_memory2_0_s2_byteenable[0]~input_o  = onchip_memory2_0_s2_byteenable[0];

assign \onchip_memory2_0_s1_writedata[1]~input_o  = onchip_memory2_0_s1_writedata[1];

assign \onchip_memory2_0_s2_writedata[1]~input_o  = onchip_memory2_0_s2_writedata[1];

assign \onchip_memory2_0_s1_writedata[2]~input_o  = onchip_memory2_0_s1_writedata[2];

assign \onchip_memory2_0_s2_writedata[2]~input_o  = onchip_memory2_0_s2_writedata[2];

assign \onchip_memory2_0_s1_writedata[3]~input_o  = onchip_memory2_0_s1_writedata[3];

assign \onchip_memory2_0_s2_writedata[3]~input_o  = onchip_memory2_0_s2_writedata[3];

assign \onchip_memory2_0_s1_writedata[4]~input_o  = onchip_memory2_0_s1_writedata[4];

assign \onchip_memory2_0_s2_writedata[4]~input_o  = onchip_memory2_0_s2_writedata[4];

assign \onchip_memory2_0_s1_writedata[5]~input_o  = onchip_memory2_0_s1_writedata[5];

assign \onchip_memory2_0_s2_writedata[5]~input_o  = onchip_memory2_0_s2_writedata[5];

assign \onchip_memory2_0_s1_writedata[6]~input_o  = onchip_memory2_0_s1_writedata[6];

assign \onchip_memory2_0_s2_writedata[6]~input_o  = onchip_memory2_0_s2_writedata[6];

assign \onchip_memory2_0_s1_writedata[7]~input_o  = onchip_memory2_0_s1_writedata[7];

assign \onchip_memory2_0_s2_writedata[7]~input_o  = onchip_memory2_0_s2_writedata[7];

assign \onchip_memory2_0_s1_writedata[8]~input_o  = onchip_memory2_0_s1_writedata[8];

assign \onchip_memory2_0_s1_byteenable[1]~input_o  = onchip_memory2_0_s1_byteenable[1];

assign \onchip_memory2_0_s2_writedata[8]~input_o  = onchip_memory2_0_s2_writedata[8];

assign \onchip_memory2_0_s2_byteenable[1]~input_o  = onchip_memory2_0_s2_byteenable[1];

assign \onchip_memory2_0_s1_writedata[9]~input_o  = onchip_memory2_0_s1_writedata[9];

assign \onchip_memory2_0_s2_writedata[9]~input_o  = onchip_memory2_0_s2_writedata[9];

assign \onchip_memory2_0_s1_writedata[10]~input_o  = onchip_memory2_0_s1_writedata[10];

assign \onchip_memory2_0_s2_writedata[10]~input_o  = onchip_memory2_0_s2_writedata[10];

assign \onchip_memory2_0_s1_writedata[11]~input_o  = onchip_memory2_0_s1_writedata[11];

assign \onchip_memory2_0_s2_writedata[11]~input_o  = onchip_memory2_0_s2_writedata[11];

assign \onchip_memory2_0_s1_writedata[12]~input_o  = onchip_memory2_0_s1_writedata[12];

assign \onchip_memory2_0_s2_writedata[12]~input_o  = onchip_memory2_0_s2_writedata[12];

assign \onchip_memory2_0_s1_writedata[13]~input_o  = onchip_memory2_0_s1_writedata[13];

assign \onchip_memory2_0_s2_writedata[13]~input_o  = onchip_memory2_0_s2_writedata[13];

assign \onchip_memory2_0_s1_writedata[14]~input_o  = onchip_memory2_0_s1_writedata[14];

assign \onchip_memory2_0_s2_writedata[14]~input_o  = onchip_memory2_0_s2_writedata[14];

assign \onchip_memory2_0_s1_writedata[15]~input_o  = onchip_memory2_0_s1_writedata[15];

assign \onchip_memory2_0_s2_writedata[15]~input_o  = onchip_memory2_0_s2_writedata[15];

assign \onchip_memory2_0_s1_writedata[16]~input_o  = onchip_memory2_0_s1_writedata[16];

assign \onchip_memory2_0_s1_byteenable[2]~input_o  = onchip_memory2_0_s1_byteenable[2];

assign \onchip_memory2_0_s2_writedata[16]~input_o  = onchip_memory2_0_s2_writedata[16];

assign \onchip_memory2_0_s2_byteenable[2]~input_o  = onchip_memory2_0_s2_byteenable[2];

assign \onchip_memory2_0_s1_writedata[17]~input_o  = onchip_memory2_0_s1_writedata[17];

assign \onchip_memory2_0_s2_writedata[17]~input_o  = onchip_memory2_0_s2_writedata[17];

assign \onchip_memory2_0_s1_writedata[18]~input_o  = onchip_memory2_0_s1_writedata[18];

assign \onchip_memory2_0_s2_writedata[18]~input_o  = onchip_memory2_0_s2_writedata[18];

assign \onchip_memory2_0_s1_writedata[19]~input_o  = onchip_memory2_0_s1_writedata[19];

assign \onchip_memory2_0_s2_writedata[19]~input_o  = onchip_memory2_0_s2_writedata[19];

assign \onchip_memory2_0_s1_writedata[20]~input_o  = onchip_memory2_0_s1_writedata[20];

assign \onchip_memory2_0_s2_writedata[20]~input_o  = onchip_memory2_0_s2_writedata[20];

assign \onchip_memory2_0_s1_writedata[21]~input_o  = onchip_memory2_0_s1_writedata[21];

assign \onchip_memory2_0_s2_writedata[21]~input_o  = onchip_memory2_0_s2_writedata[21];

assign \onchip_memory2_0_s1_writedata[22]~input_o  = onchip_memory2_0_s1_writedata[22];

assign \onchip_memory2_0_s2_writedata[22]~input_o  = onchip_memory2_0_s2_writedata[22];

assign \onchip_memory2_0_s1_writedata[23]~input_o  = onchip_memory2_0_s1_writedata[23];

assign \onchip_memory2_0_s2_writedata[23]~input_o  = onchip_memory2_0_s2_writedata[23];

assign \onchip_memory2_0_s1_writedata[24]~input_o  = onchip_memory2_0_s1_writedata[24];

assign \onchip_memory2_0_s1_byteenable[3]~input_o  = onchip_memory2_0_s1_byteenable[3];

assign \onchip_memory2_0_s2_writedata[24]~input_o  = onchip_memory2_0_s2_writedata[24];

assign \onchip_memory2_0_s2_byteenable[3]~input_o  = onchip_memory2_0_s2_byteenable[3];

assign \onchip_memory2_0_s1_writedata[25]~input_o  = onchip_memory2_0_s1_writedata[25];

assign \onchip_memory2_0_s2_writedata[25]~input_o  = onchip_memory2_0_s2_writedata[25];

assign \onchip_memory2_0_s1_writedata[26]~input_o  = onchip_memory2_0_s1_writedata[26];

assign \onchip_memory2_0_s2_writedata[26]~input_o  = onchip_memory2_0_s2_writedata[26];

assign \onchip_memory2_0_s1_writedata[27]~input_o  = onchip_memory2_0_s1_writedata[27];

assign \onchip_memory2_0_s2_writedata[27]~input_o  = onchip_memory2_0_s2_writedata[27];

assign \onchip_memory2_0_s1_writedata[28]~input_o  = onchip_memory2_0_s1_writedata[28];

assign \onchip_memory2_0_s2_writedata[28]~input_o  = onchip_memory2_0_s2_writedata[28];

assign \onchip_memory2_0_s1_writedata[29]~input_o  = onchip_memory2_0_s1_writedata[29];

assign \onchip_memory2_0_s2_writedata[29]~input_o  = onchip_memory2_0_s2_writedata[29];

assign \onchip_memory2_0_s1_writedata[30]~input_o  = onchip_memory2_0_s1_writedata[30];

assign \onchip_memory2_0_s2_writedata[30]~input_o  = onchip_memory2_0_s2_writedata[30];

assign \onchip_memory2_0_s1_writedata[31]~input_o  = onchip_memory2_0_s1_writedata[31];

assign \onchip_memory2_0_s2_writedata[31]~input_o  = onchip_memory2_0_s2_writedata[31];

assign \onchip_memory2_0_s1_writedata[32]~input_o  = onchip_memory2_0_s1_writedata[32];

assign \onchip_memory2_0_s1_byteenable[4]~input_o  = onchip_memory2_0_s1_byteenable[4];

assign \onchip_memory2_0_s2_writedata[32]~input_o  = onchip_memory2_0_s2_writedata[32];

assign \onchip_memory2_0_s2_byteenable[4]~input_o  = onchip_memory2_0_s2_byteenable[4];

assign \onchip_memory2_0_s1_writedata[33]~input_o  = onchip_memory2_0_s1_writedata[33];

assign \onchip_memory2_0_s2_writedata[33]~input_o  = onchip_memory2_0_s2_writedata[33];

assign \onchip_memory2_0_s1_writedata[34]~input_o  = onchip_memory2_0_s1_writedata[34];

assign \onchip_memory2_0_s2_writedata[34]~input_o  = onchip_memory2_0_s2_writedata[34];

assign \onchip_memory2_0_s1_writedata[35]~input_o  = onchip_memory2_0_s1_writedata[35];

assign \onchip_memory2_0_s2_writedata[35]~input_o  = onchip_memory2_0_s2_writedata[35];

assign \onchip_memory2_0_s1_writedata[36]~input_o  = onchip_memory2_0_s1_writedata[36];

assign \onchip_memory2_0_s2_writedata[36]~input_o  = onchip_memory2_0_s2_writedata[36];

assign \onchip_memory2_0_s1_writedata[37]~input_o  = onchip_memory2_0_s1_writedata[37];

assign \onchip_memory2_0_s2_writedata[37]~input_o  = onchip_memory2_0_s2_writedata[37];

assign \onchip_memory2_0_s1_writedata[38]~input_o  = onchip_memory2_0_s1_writedata[38];

assign \onchip_memory2_0_s2_writedata[38]~input_o  = onchip_memory2_0_s2_writedata[38];

assign \onchip_memory2_0_s1_writedata[39]~input_o  = onchip_memory2_0_s1_writedata[39];

assign \onchip_memory2_0_s2_writedata[39]~input_o  = onchip_memory2_0_s2_writedata[39];

assign \onchip_memory2_0_s1_writedata[40]~input_o  = onchip_memory2_0_s1_writedata[40];

assign \onchip_memory2_0_s1_byteenable[5]~input_o  = onchip_memory2_0_s1_byteenable[5];

assign \onchip_memory2_0_s2_writedata[40]~input_o  = onchip_memory2_0_s2_writedata[40];

assign \onchip_memory2_0_s2_byteenable[5]~input_o  = onchip_memory2_0_s2_byteenable[5];

assign \onchip_memory2_0_s1_writedata[41]~input_o  = onchip_memory2_0_s1_writedata[41];

assign \onchip_memory2_0_s2_writedata[41]~input_o  = onchip_memory2_0_s2_writedata[41];

assign \onchip_memory2_0_s1_writedata[42]~input_o  = onchip_memory2_0_s1_writedata[42];

assign \onchip_memory2_0_s2_writedata[42]~input_o  = onchip_memory2_0_s2_writedata[42];

assign \onchip_memory2_0_s1_writedata[43]~input_o  = onchip_memory2_0_s1_writedata[43];

assign \onchip_memory2_0_s2_writedata[43]~input_o  = onchip_memory2_0_s2_writedata[43];

assign \onchip_memory2_0_s1_writedata[44]~input_o  = onchip_memory2_0_s1_writedata[44];

assign \onchip_memory2_0_s2_writedata[44]~input_o  = onchip_memory2_0_s2_writedata[44];

assign \onchip_memory2_0_s1_writedata[45]~input_o  = onchip_memory2_0_s1_writedata[45];

assign \onchip_memory2_0_s2_writedata[45]~input_o  = onchip_memory2_0_s2_writedata[45];

assign \onchip_memory2_0_s1_writedata[46]~input_o  = onchip_memory2_0_s1_writedata[46];

assign \onchip_memory2_0_s2_writedata[46]~input_o  = onchip_memory2_0_s2_writedata[46];

assign \onchip_memory2_0_s1_writedata[47]~input_o  = onchip_memory2_0_s1_writedata[47];

assign \onchip_memory2_0_s2_writedata[47]~input_o  = onchip_memory2_0_s2_writedata[47];

assign \onchip_memory2_0_s1_writedata[48]~input_o  = onchip_memory2_0_s1_writedata[48];

assign \onchip_memory2_0_s1_byteenable[6]~input_o  = onchip_memory2_0_s1_byteenable[6];

assign \onchip_memory2_0_s2_writedata[48]~input_o  = onchip_memory2_0_s2_writedata[48];

assign \onchip_memory2_0_s2_byteenable[6]~input_o  = onchip_memory2_0_s2_byteenable[6];

assign \onchip_memory2_0_s1_writedata[49]~input_o  = onchip_memory2_0_s1_writedata[49];

assign \onchip_memory2_0_s2_writedata[49]~input_o  = onchip_memory2_0_s2_writedata[49];

assign \onchip_memory2_0_s1_writedata[50]~input_o  = onchip_memory2_0_s1_writedata[50];

assign \onchip_memory2_0_s2_writedata[50]~input_o  = onchip_memory2_0_s2_writedata[50];

assign \onchip_memory2_0_s1_writedata[51]~input_o  = onchip_memory2_0_s1_writedata[51];

assign \onchip_memory2_0_s2_writedata[51]~input_o  = onchip_memory2_0_s2_writedata[51];

assign \onchip_memory2_0_s1_writedata[52]~input_o  = onchip_memory2_0_s1_writedata[52];

assign \onchip_memory2_0_s2_writedata[52]~input_o  = onchip_memory2_0_s2_writedata[52];

assign \onchip_memory2_0_s1_writedata[53]~input_o  = onchip_memory2_0_s1_writedata[53];

assign \onchip_memory2_0_s2_writedata[53]~input_o  = onchip_memory2_0_s2_writedata[53];

assign \onchip_memory2_0_s1_writedata[54]~input_o  = onchip_memory2_0_s1_writedata[54];

assign \onchip_memory2_0_s2_writedata[54]~input_o  = onchip_memory2_0_s2_writedata[54];

assign \onchip_memory2_0_s1_writedata[55]~input_o  = onchip_memory2_0_s1_writedata[55];

assign \onchip_memory2_0_s2_writedata[55]~input_o  = onchip_memory2_0_s2_writedata[55];

assign \onchip_memory2_0_s1_writedata[56]~input_o  = onchip_memory2_0_s1_writedata[56];

assign \onchip_memory2_0_s1_byteenable[7]~input_o  = onchip_memory2_0_s1_byteenable[7];

assign \onchip_memory2_0_s2_writedata[56]~input_o  = onchip_memory2_0_s2_writedata[56];

assign \onchip_memory2_0_s2_byteenable[7]~input_o  = onchip_memory2_0_s2_byteenable[7];

assign \onchip_memory2_0_s1_writedata[57]~input_o  = onchip_memory2_0_s1_writedata[57];

assign \onchip_memory2_0_s2_writedata[57]~input_o  = onchip_memory2_0_s2_writedata[57];

assign \onchip_memory2_0_s1_writedata[58]~input_o  = onchip_memory2_0_s1_writedata[58];

assign \onchip_memory2_0_s2_writedata[58]~input_o  = onchip_memory2_0_s2_writedata[58];

assign \onchip_memory2_0_s1_writedata[59]~input_o  = onchip_memory2_0_s1_writedata[59];

assign \onchip_memory2_0_s2_writedata[59]~input_o  = onchip_memory2_0_s2_writedata[59];

assign \onchip_memory2_0_s1_writedata[60]~input_o  = onchip_memory2_0_s1_writedata[60];

assign \onchip_memory2_0_s2_writedata[60]~input_o  = onchip_memory2_0_s2_writedata[60];

assign \onchip_memory2_0_s1_writedata[61]~input_o  = onchip_memory2_0_s1_writedata[61];

assign \onchip_memory2_0_s2_writedata[61]~input_o  = onchip_memory2_0_s2_writedata[61];

assign \onchip_memory2_0_s1_writedata[62]~input_o  = onchip_memory2_0_s1_writedata[62];

assign \onchip_memory2_0_s2_writedata[62]~input_o  = onchip_memory2_0_s2_writedata[62];

assign \onchip_memory2_0_s1_writedata[63]~input_o  = onchip_memory2_0_s1_writedata[63];

assign \onchip_memory2_0_s2_writedata[63]~input_o  = onchip_memory2_0_s2_writedata[63];

assign \reset_reset_n~input_o  = reset_reset_n;

assign onchip_memory2_0_s1_readdata[0] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[0]~0_combout ;

assign onchip_memory2_0_s1_readdata[1] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[1]~1_combout ;

assign onchip_memory2_0_s1_readdata[2] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[2]~2_combout ;

assign onchip_memory2_0_s1_readdata[3] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[3]~3_combout ;

assign onchip_memory2_0_s1_readdata[4] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[4]~4_combout ;

assign onchip_memory2_0_s1_readdata[5] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[5]~5_combout ;

assign onchip_memory2_0_s1_readdata[6] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[6]~6_combout ;

assign onchip_memory2_0_s1_readdata[7] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[7]~7_combout ;

assign onchip_memory2_0_s1_readdata[8] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[8]~8_combout ;

assign onchip_memory2_0_s1_readdata[9] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[9]~9_combout ;

assign onchip_memory2_0_s1_readdata[10] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[10]~10_combout ;

assign onchip_memory2_0_s1_readdata[11] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[11]~11_combout ;

assign onchip_memory2_0_s1_readdata[12] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[12]~12_combout ;

assign onchip_memory2_0_s1_readdata[13] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[13]~13_combout ;

assign onchip_memory2_0_s1_readdata[14] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[14]~14_combout ;

assign onchip_memory2_0_s1_readdata[15] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[15]~15_combout ;

assign onchip_memory2_0_s1_readdata[16] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[16]~16_combout ;

assign onchip_memory2_0_s1_readdata[17] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[17]~17_combout ;

assign onchip_memory2_0_s1_readdata[18] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[18]~18_combout ;

assign onchip_memory2_0_s1_readdata[19] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[19]~19_combout ;

assign onchip_memory2_0_s1_readdata[20] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[20]~20_combout ;

assign onchip_memory2_0_s1_readdata[21] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[21]~21_combout ;

assign onchip_memory2_0_s1_readdata[22] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[22]~22_combout ;

assign onchip_memory2_0_s1_readdata[23] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[23]~23_combout ;

assign onchip_memory2_0_s1_readdata[24] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[24]~24_combout ;

assign onchip_memory2_0_s1_readdata[25] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[25]~25_combout ;

assign onchip_memory2_0_s1_readdata[26] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[26]~26_combout ;

assign onchip_memory2_0_s1_readdata[27] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[27]~27_combout ;

assign onchip_memory2_0_s1_readdata[28] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[28]~28_combout ;

assign onchip_memory2_0_s1_readdata[29] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[29]~29_combout ;

assign onchip_memory2_0_s1_readdata[30] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[30]~30_combout ;

assign onchip_memory2_0_s1_readdata[31] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[31]~31_combout ;

assign onchip_memory2_0_s1_readdata[32] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[32]~32_combout ;

assign onchip_memory2_0_s1_readdata[33] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[33]~33_combout ;

assign onchip_memory2_0_s1_readdata[34] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[34]~34_combout ;

assign onchip_memory2_0_s1_readdata[35] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[35]~35_combout ;

assign onchip_memory2_0_s1_readdata[36] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[36]~36_combout ;

assign onchip_memory2_0_s1_readdata[37] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[37]~37_combout ;

assign onchip_memory2_0_s1_readdata[38] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[38]~38_combout ;

assign onchip_memory2_0_s1_readdata[39] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[39]~39_combout ;

assign onchip_memory2_0_s1_readdata[40] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[40]~40_combout ;

assign onchip_memory2_0_s1_readdata[41] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[41]~41_combout ;

assign onchip_memory2_0_s1_readdata[42] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[42]~42_combout ;

assign onchip_memory2_0_s1_readdata[43] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[43]~43_combout ;

assign onchip_memory2_0_s1_readdata[44] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[44]~44_combout ;

assign onchip_memory2_0_s1_readdata[45] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[45]~45_combout ;

assign onchip_memory2_0_s1_readdata[46] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[46]~46_combout ;

assign onchip_memory2_0_s1_readdata[47] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[47]~47_combout ;

assign onchip_memory2_0_s1_readdata[48] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[48]~48_combout ;

assign onchip_memory2_0_s1_readdata[49] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[49]~49_combout ;

assign onchip_memory2_0_s1_readdata[50] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[50]~50_combout ;

assign onchip_memory2_0_s1_readdata[51] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[51]~51_combout ;

assign onchip_memory2_0_s1_readdata[52] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[52]~52_combout ;

assign onchip_memory2_0_s1_readdata[53] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[53]~53_combout ;

assign onchip_memory2_0_s1_readdata[54] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[54]~54_combout ;

assign onchip_memory2_0_s1_readdata[55] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[55]~55_combout ;

assign onchip_memory2_0_s1_readdata[56] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[56]~56_combout ;

assign onchip_memory2_0_s1_readdata[57] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[57]~57_combout ;

assign onchip_memory2_0_s1_readdata[58] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[58]~58_combout ;

assign onchip_memory2_0_s1_readdata[59] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[59]~59_combout ;

assign onchip_memory2_0_s1_readdata[60] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[60]~60_combout ;

assign onchip_memory2_0_s1_readdata[61] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[61]~61_combout ;

assign onchip_memory2_0_s1_readdata[62] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[62]~62_combout ;

assign onchip_memory2_0_s1_readdata[63] = \onchip_memory2_0|the_altsyncram|auto_generated|mux4|result_node[63]~63_combout ;

assign onchip_memory2_0_s2_readdata[0] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[0]~0_combout ;

assign onchip_memory2_0_s2_readdata[1] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[1]~1_combout ;

assign onchip_memory2_0_s2_readdata[2] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[2]~2_combout ;

assign onchip_memory2_0_s2_readdata[3] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[3]~3_combout ;

assign onchip_memory2_0_s2_readdata[4] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[4]~4_combout ;

assign onchip_memory2_0_s2_readdata[5] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[5]~5_combout ;

assign onchip_memory2_0_s2_readdata[6] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[6]~6_combout ;

assign onchip_memory2_0_s2_readdata[7] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[7]~7_combout ;

assign onchip_memory2_0_s2_readdata[8] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[8]~8_combout ;

assign onchip_memory2_0_s2_readdata[9] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[9]~9_combout ;

assign onchip_memory2_0_s2_readdata[10] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[10]~10_combout ;

assign onchip_memory2_0_s2_readdata[11] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[11]~11_combout ;

assign onchip_memory2_0_s2_readdata[12] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[12]~12_combout ;

assign onchip_memory2_0_s2_readdata[13] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[13]~13_combout ;

assign onchip_memory2_0_s2_readdata[14] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[14]~14_combout ;

assign onchip_memory2_0_s2_readdata[15] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[15]~15_combout ;

assign onchip_memory2_0_s2_readdata[16] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[16]~16_combout ;

assign onchip_memory2_0_s2_readdata[17] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[17]~17_combout ;

assign onchip_memory2_0_s2_readdata[18] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[18]~18_combout ;

assign onchip_memory2_0_s2_readdata[19] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[19]~19_combout ;

assign onchip_memory2_0_s2_readdata[20] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[20]~20_combout ;

assign onchip_memory2_0_s2_readdata[21] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[21]~21_combout ;

assign onchip_memory2_0_s2_readdata[22] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[22]~22_combout ;

assign onchip_memory2_0_s2_readdata[23] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[23]~23_combout ;

assign onchip_memory2_0_s2_readdata[24] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[24]~24_combout ;

assign onchip_memory2_0_s2_readdata[25] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[25]~25_combout ;

assign onchip_memory2_0_s2_readdata[26] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[26]~26_combout ;

assign onchip_memory2_0_s2_readdata[27] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[27]~27_combout ;

assign onchip_memory2_0_s2_readdata[28] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[28]~28_combout ;

assign onchip_memory2_0_s2_readdata[29] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[29]~29_combout ;

assign onchip_memory2_0_s2_readdata[30] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[30]~30_combout ;

assign onchip_memory2_0_s2_readdata[31] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[31]~31_combout ;

assign onchip_memory2_0_s2_readdata[32] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[32]~32_combout ;

assign onchip_memory2_0_s2_readdata[33] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[33]~33_combout ;

assign onchip_memory2_0_s2_readdata[34] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[34]~34_combout ;

assign onchip_memory2_0_s2_readdata[35] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[35]~35_combout ;

assign onchip_memory2_0_s2_readdata[36] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[36]~36_combout ;

assign onchip_memory2_0_s2_readdata[37] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[37]~37_combout ;

assign onchip_memory2_0_s2_readdata[38] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[38]~38_combout ;

assign onchip_memory2_0_s2_readdata[39] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[39]~39_combout ;

assign onchip_memory2_0_s2_readdata[40] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[40]~40_combout ;

assign onchip_memory2_0_s2_readdata[41] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[41]~41_combout ;

assign onchip_memory2_0_s2_readdata[42] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[42]~42_combout ;

assign onchip_memory2_0_s2_readdata[43] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[43]~43_combout ;

assign onchip_memory2_0_s2_readdata[44] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[44]~44_combout ;

assign onchip_memory2_0_s2_readdata[45] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[45]~45_combout ;

assign onchip_memory2_0_s2_readdata[46] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[46]~46_combout ;

assign onchip_memory2_0_s2_readdata[47] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[47]~47_combout ;

assign onchip_memory2_0_s2_readdata[48] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[48]~48_combout ;

assign onchip_memory2_0_s2_readdata[49] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[49]~49_combout ;

assign onchip_memory2_0_s2_readdata[50] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[50]~50_combout ;

assign onchip_memory2_0_s2_readdata[51] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[51]~51_combout ;

assign onchip_memory2_0_s2_readdata[52] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[52]~52_combout ;

assign onchip_memory2_0_s2_readdata[53] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[53]~53_combout ;

assign onchip_memory2_0_s2_readdata[54] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[54]~54_combout ;

assign onchip_memory2_0_s2_readdata[55] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[55]~55_combout ;

assign onchip_memory2_0_s2_readdata[56] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[56]~56_combout ;

assign onchip_memory2_0_s2_readdata[57] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[57]~57_combout ;

assign onchip_memory2_0_s2_readdata[58] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[58]~58_combout ;

assign onchip_memory2_0_s2_readdata[59] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[59]~59_combout ;

assign onchip_memory2_0_s2_readdata[60] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[60]~60_combout ;

assign onchip_memory2_0_s2_readdata[61] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[61]~61_combout ;

assign onchip_memory2_0_s2_readdata[62] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[62]~62_combout ;

assign onchip_memory2_0_s2_readdata[63] = \onchip_memory2_0|the_altsyncram|auto_generated|mux5|result_node[63]~63_combout ;

endmodule

module qtestpd_altera_reset_controller (
	r_early_rst1,
	clk_clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	r_early_rst1;
input 	clk_clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \always2~0_combout ;


qtestpd_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk));

qtestpd_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.clk(clk_clk),
	.reset_reset_n(reset_reset_n));

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cycloneiv_lcell_comb \r_sync_rst_chain~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_reset_synchronizer_int_chain[2]~q ),
	.datad(\r_sync_rst_chain[3]~q ),
	.cin(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.cout());
defparam \r_sync_rst_chain~0 .lut_mask = 16'hF000;
defparam \r_sync_rst_chain~0 .sum_lutc_input = "datac";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cycloneiv_lcell_comb \always2~0 (
	.dataa(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\r_sync_rst_chain[2]~q ),
	.cin(gnd),
	.combout(\always2~0_combout ),
	.cout());
defparam \always2~0 .lut_mask = 16'hAAFF;
defparam \always2~0 .sum_lutc_input = "datac";

endmodule

module qtestpd_altera_reset_synchronizer (
	altera_reset_synchronizer_int_chain_out1,
	clk)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cycloneiv_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.cout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 16'h0000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .sum_lutc_input = "datac";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module qtestpd_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	clk,
	reset_reset_n)/* synthesis synthesis_greybox=0 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	clk;
input 	reset_reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(reset_reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module qtestpd_qtestpd_onchip_memory2_0 (
	result_node_0,
	result_node_1,
	result_node_2,
	result_node_3,
	result_node_4,
	result_node_5,
	result_node_6,
	result_node_7,
	result_node_8,
	result_node_9,
	result_node_10,
	result_node_11,
	result_node_12,
	result_node_13,
	result_node_14,
	result_node_15,
	result_node_16,
	result_node_17,
	result_node_18,
	result_node_19,
	result_node_20,
	result_node_21,
	result_node_22,
	result_node_23,
	result_node_24,
	result_node_25,
	result_node_26,
	result_node_27,
	result_node_28,
	result_node_29,
	result_node_30,
	result_node_31,
	result_node_32,
	result_node_33,
	result_node_34,
	result_node_35,
	result_node_36,
	result_node_37,
	result_node_38,
	result_node_39,
	result_node_40,
	result_node_41,
	result_node_42,
	result_node_43,
	result_node_44,
	result_node_45,
	result_node_46,
	result_node_47,
	result_node_48,
	result_node_49,
	result_node_50,
	result_node_51,
	result_node_52,
	result_node_53,
	result_node_54,
	result_node_55,
	result_node_56,
	result_node_57,
	result_node_58,
	result_node_59,
	result_node_60,
	result_node_61,
	result_node_62,
	result_node_63,
	result_node_01,
	result_node_110,
	result_node_210,
	result_node_310,
	result_node_410,
	result_node_510,
	result_node_64,
	result_node_71,
	result_node_81,
	result_node_91,
	result_node_101,
	result_node_111,
	result_node_121,
	result_node_131,
	result_node_141,
	result_node_151,
	result_node_161,
	result_node_171,
	result_node_181,
	result_node_191,
	result_node_201,
	result_node_211,
	result_node_221,
	result_node_231,
	result_node_241,
	result_node_251,
	result_node_261,
	result_node_271,
	result_node_281,
	result_node_291,
	result_node_301,
	result_node_311,
	result_node_321,
	result_node_331,
	result_node_341,
	result_node_351,
	result_node_361,
	result_node_371,
	result_node_381,
	result_node_391,
	result_node_401,
	result_node_411,
	result_node_421,
	result_node_431,
	result_node_441,
	result_node_451,
	result_node_461,
	result_node_471,
	result_node_481,
	result_node_491,
	result_node_501,
	result_node_511,
	result_node_521,
	result_node_531,
	result_node_541,
	result_node_551,
	result_node_561,
	result_node_571,
	result_node_581,
	result_node_591,
	result_node_601,
	result_node_611,
	result_node_621,
	result_node_631,
	r_early_rst,
	onchip_memory2_0_s1_address_13,
	onchip_memory2_0_s1_chipselect,
	onchip_memory2_0_s1_write,
	onchip_memory2_0_s2_address_13,
	onchip_memory2_0_s2_chipselect,
	onchip_memory2_0_s2_write,
	clk_clk,
	onchip_memory2_0_s1_clken,
	onchip_memory2_0_s2_clken,
	onchip_memory2_0_s1_writedata_0,
	onchip_memory2_0_s1_address_0,
	onchip_memory2_0_s1_address_1,
	onchip_memory2_0_s1_address_2,
	onchip_memory2_0_s1_address_3,
	onchip_memory2_0_s1_address_4,
	onchip_memory2_0_s1_address_5,
	onchip_memory2_0_s1_address_6,
	onchip_memory2_0_s1_address_7,
	onchip_memory2_0_s1_address_8,
	onchip_memory2_0_s1_address_9,
	onchip_memory2_0_s1_address_10,
	onchip_memory2_0_s1_address_11,
	onchip_memory2_0_s1_address_12,
	onchip_memory2_0_s1_byteenable_0,
	onchip_memory2_0_s2_writedata_0,
	onchip_memory2_0_s2_address_0,
	onchip_memory2_0_s2_address_1,
	onchip_memory2_0_s2_address_2,
	onchip_memory2_0_s2_address_3,
	onchip_memory2_0_s2_address_4,
	onchip_memory2_0_s2_address_5,
	onchip_memory2_0_s2_address_6,
	onchip_memory2_0_s2_address_7,
	onchip_memory2_0_s2_address_8,
	onchip_memory2_0_s2_address_9,
	onchip_memory2_0_s2_address_10,
	onchip_memory2_0_s2_address_11,
	onchip_memory2_0_s2_address_12,
	onchip_memory2_0_s2_byteenable_0,
	onchip_memory2_0_s1_writedata_1,
	onchip_memory2_0_s2_writedata_1,
	onchip_memory2_0_s1_writedata_2,
	onchip_memory2_0_s2_writedata_2,
	onchip_memory2_0_s1_writedata_3,
	onchip_memory2_0_s2_writedata_3,
	onchip_memory2_0_s1_writedata_4,
	onchip_memory2_0_s2_writedata_4,
	onchip_memory2_0_s1_writedata_5,
	onchip_memory2_0_s2_writedata_5,
	onchip_memory2_0_s1_writedata_6,
	onchip_memory2_0_s2_writedata_6,
	onchip_memory2_0_s1_writedata_7,
	onchip_memory2_0_s2_writedata_7,
	onchip_memory2_0_s1_writedata_8,
	onchip_memory2_0_s1_byteenable_1,
	onchip_memory2_0_s2_writedata_8,
	onchip_memory2_0_s2_byteenable_1,
	onchip_memory2_0_s1_writedata_9,
	onchip_memory2_0_s2_writedata_9,
	onchip_memory2_0_s1_writedata_10,
	onchip_memory2_0_s2_writedata_10,
	onchip_memory2_0_s1_writedata_11,
	onchip_memory2_0_s2_writedata_11,
	onchip_memory2_0_s1_writedata_12,
	onchip_memory2_0_s2_writedata_12,
	onchip_memory2_0_s1_writedata_13,
	onchip_memory2_0_s2_writedata_13,
	onchip_memory2_0_s1_writedata_14,
	onchip_memory2_0_s2_writedata_14,
	onchip_memory2_0_s1_writedata_15,
	onchip_memory2_0_s2_writedata_15,
	onchip_memory2_0_s1_writedata_16,
	onchip_memory2_0_s1_byteenable_2,
	onchip_memory2_0_s2_writedata_16,
	onchip_memory2_0_s2_byteenable_2,
	onchip_memory2_0_s1_writedata_17,
	onchip_memory2_0_s2_writedata_17,
	onchip_memory2_0_s1_writedata_18,
	onchip_memory2_0_s2_writedata_18,
	onchip_memory2_0_s1_writedata_19,
	onchip_memory2_0_s2_writedata_19,
	onchip_memory2_0_s1_writedata_20,
	onchip_memory2_0_s2_writedata_20,
	onchip_memory2_0_s1_writedata_21,
	onchip_memory2_0_s2_writedata_21,
	onchip_memory2_0_s1_writedata_22,
	onchip_memory2_0_s2_writedata_22,
	onchip_memory2_0_s1_writedata_23,
	onchip_memory2_0_s2_writedata_23,
	onchip_memory2_0_s1_writedata_24,
	onchip_memory2_0_s1_byteenable_3,
	onchip_memory2_0_s2_writedata_24,
	onchip_memory2_0_s2_byteenable_3,
	onchip_memory2_0_s1_writedata_25,
	onchip_memory2_0_s2_writedata_25,
	onchip_memory2_0_s1_writedata_26,
	onchip_memory2_0_s2_writedata_26,
	onchip_memory2_0_s1_writedata_27,
	onchip_memory2_0_s2_writedata_27,
	onchip_memory2_0_s1_writedata_28,
	onchip_memory2_0_s2_writedata_28,
	onchip_memory2_0_s1_writedata_29,
	onchip_memory2_0_s2_writedata_29,
	onchip_memory2_0_s1_writedata_30,
	onchip_memory2_0_s2_writedata_30,
	onchip_memory2_0_s1_writedata_31,
	onchip_memory2_0_s2_writedata_31,
	onchip_memory2_0_s1_writedata_32,
	onchip_memory2_0_s1_byteenable_4,
	onchip_memory2_0_s2_writedata_32,
	onchip_memory2_0_s2_byteenable_4,
	onchip_memory2_0_s1_writedata_33,
	onchip_memory2_0_s2_writedata_33,
	onchip_memory2_0_s1_writedata_34,
	onchip_memory2_0_s2_writedata_34,
	onchip_memory2_0_s1_writedata_35,
	onchip_memory2_0_s2_writedata_35,
	onchip_memory2_0_s1_writedata_36,
	onchip_memory2_0_s2_writedata_36,
	onchip_memory2_0_s1_writedata_37,
	onchip_memory2_0_s2_writedata_37,
	onchip_memory2_0_s1_writedata_38,
	onchip_memory2_0_s2_writedata_38,
	onchip_memory2_0_s1_writedata_39,
	onchip_memory2_0_s2_writedata_39,
	onchip_memory2_0_s1_writedata_40,
	onchip_memory2_0_s1_byteenable_5,
	onchip_memory2_0_s2_writedata_40,
	onchip_memory2_0_s2_byteenable_5,
	onchip_memory2_0_s1_writedata_41,
	onchip_memory2_0_s2_writedata_41,
	onchip_memory2_0_s1_writedata_42,
	onchip_memory2_0_s2_writedata_42,
	onchip_memory2_0_s1_writedata_43,
	onchip_memory2_0_s2_writedata_43,
	onchip_memory2_0_s1_writedata_44,
	onchip_memory2_0_s2_writedata_44,
	onchip_memory2_0_s1_writedata_45,
	onchip_memory2_0_s2_writedata_45,
	onchip_memory2_0_s1_writedata_46,
	onchip_memory2_0_s2_writedata_46,
	onchip_memory2_0_s1_writedata_47,
	onchip_memory2_0_s2_writedata_47,
	onchip_memory2_0_s1_writedata_48,
	onchip_memory2_0_s1_byteenable_6,
	onchip_memory2_0_s2_writedata_48,
	onchip_memory2_0_s2_byteenable_6,
	onchip_memory2_0_s1_writedata_49,
	onchip_memory2_0_s2_writedata_49,
	onchip_memory2_0_s1_writedata_50,
	onchip_memory2_0_s2_writedata_50,
	onchip_memory2_0_s1_writedata_51,
	onchip_memory2_0_s2_writedata_51,
	onchip_memory2_0_s1_writedata_52,
	onchip_memory2_0_s2_writedata_52,
	onchip_memory2_0_s1_writedata_53,
	onchip_memory2_0_s2_writedata_53,
	onchip_memory2_0_s1_writedata_54,
	onchip_memory2_0_s2_writedata_54,
	onchip_memory2_0_s1_writedata_55,
	onchip_memory2_0_s2_writedata_55,
	onchip_memory2_0_s1_writedata_56,
	onchip_memory2_0_s1_byteenable_7,
	onchip_memory2_0_s2_writedata_56,
	onchip_memory2_0_s2_byteenable_7,
	onchip_memory2_0_s1_writedata_57,
	onchip_memory2_0_s2_writedata_57,
	onchip_memory2_0_s1_writedata_58,
	onchip_memory2_0_s2_writedata_58,
	onchip_memory2_0_s1_writedata_59,
	onchip_memory2_0_s2_writedata_59,
	onchip_memory2_0_s1_writedata_60,
	onchip_memory2_0_s2_writedata_60,
	onchip_memory2_0_s1_writedata_61,
	onchip_memory2_0_s2_writedata_61,
	onchip_memory2_0_s1_writedata_62,
	onchip_memory2_0_s2_writedata_62,
	onchip_memory2_0_s1_writedata_63,
	onchip_memory2_0_s2_writedata_63)/* synthesis synthesis_greybox=0 */;
output 	result_node_0;
output 	result_node_1;
output 	result_node_2;
output 	result_node_3;
output 	result_node_4;
output 	result_node_5;
output 	result_node_6;
output 	result_node_7;
output 	result_node_8;
output 	result_node_9;
output 	result_node_10;
output 	result_node_11;
output 	result_node_12;
output 	result_node_13;
output 	result_node_14;
output 	result_node_15;
output 	result_node_16;
output 	result_node_17;
output 	result_node_18;
output 	result_node_19;
output 	result_node_20;
output 	result_node_21;
output 	result_node_22;
output 	result_node_23;
output 	result_node_24;
output 	result_node_25;
output 	result_node_26;
output 	result_node_27;
output 	result_node_28;
output 	result_node_29;
output 	result_node_30;
output 	result_node_31;
output 	result_node_32;
output 	result_node_33;
output 	result_node_34;
output 	result_node_35;
output 	result_node_36;
output 	result_node_37;
output 	result_node_38;
output 	result_node_39;
output 	result_node_40;
output 	result_node_41;
output 	result_node_42;
output 	result_node_43;
output 	result_node_44;
output 	result_node_45;
output 	result_node_46;
output 	result_node_47;
output 	result_node_48;
output 	result_node_49;
output 	result_node_50;
output 	result_node_51;
output 	result_node_52;
output 	result_node_53;
output 	result_node_54;
output 	result_node_55;
output 	result_node_56;
output 	result_node_57;
output 	result_node_58;
output 	result_node_59;
output 	result_node_60;
output 	result_node_61;
output 	result_node_62;
output 	result_node_63;
output 	result_node_01;
output 	result_node_110;
output 	result_node_210;
output 	result_node_310;
output 	result_node_410;
output 	result_node_510;
output 	result_node_64;
output 	result_node_71;
output 	result_node_81;
output 	result_node_91;
output 	result_node_101;
output 	result_node_111;
output 	result_node_121;
output 	result_node_131;
output 	result_node_141;
output 	result_node_151;
output 	result_node_161;
output 	result_node_171;
output 	result_node_181;
output 	result_node_191;
output 	result_node_201;
output 	result_node_211;
output 	result_node_221;
output 	result_node_231;
output 	result_node_241;
output 	result_node_251;
output 	result_node_261;
output 	result_node_271;
output 	result_node_281;
output 	result_node_291;
output 	result_node_301;
output 	result_node_311;
output 	result_node_321;
output 	result_node_331;
output 	result_node_341;
output 	result_node_351;
output 	result_node_361;
output 	result_node_371;
output 	result_node_381;
output 	result_node_391;
output 	result_node_401;
output 	result_node_411;
output 	result_node_421;
output 	result_node_431;
output 	result_node_441;
output 	result_node_451;
output 	result_node_461;
output 	result_node_471;
output 	result_node_481;
output 	result_node_491;
output 	result_node_501;
output 	result_node_511;
output 	result_node_521;
output 	result_node_531;
output 	result_node_541;
output 	result_node_551;
output 	result_node_561;
output 	result_node_571;
output 	result_node_581;
output 	result_node_591;
output 	result_node_601;
output 	result_node_611;
output 	result_node_621;
output 	result_node_631;
input 	r_early_rst;
input 	onchip_memory2_0_s1_address_13;
input 	onchip_memory2_0_s1_chipselect;
input 	onchip_memory2_0_s1_write;
input 	onchip_memory2_0_s2_address_13;
input 	onchip_memory2_0_s2_chipselect;
input 	onchip_memory2_0_s2_write;
input 	clk_clk;
input 	onchip_memory2_0_s1_clken;
input 	onchip_memory2_0_s2_clken;
input 	onchip_memory2_0_s1_writedata_0;
input 	onchip_memory2_0_s1_address_0;
input 	onchip_memory2_0_s1_address_1;
input 	onchip_memory2_0_s1_address_2;
input 	onchip_memory2_0_s1_address_3;
input 	onchip_memory2_0_s1_address_4;
input 	onchip_memory2_0_s1_address_5;
input 	onchip_memory2_0_s1_address_6;
input 	onchip_memory2_0_s1_address_7;
input 	onchip_memory2_0_s1_address_8;
input 	onchip_memory2_0_s1_address_9;
input 	onchip_memory2_0_s1_address_10;
input 	onchip_memory2_0_s1_address_11;
input 	onchip_memory2_0_s1_address_12;
input 	onchip_memory2_0_s1_byteenable_0;
input 	onchip_memory2_0_s2_writedata_0;
input 	onchip_memory2_0_s2_address_0;
input 	onchip_memory2_0_s2_address_1;
input 	onchip_memory2_0_s2_address_2;
input 	onchip_memory2_0_s2_address_3;
input 	onchip_memory2_0_s2_address_4;
input 	onchip_memory2_0_s2_address_5;
input 	onchip_memory2_0_s2_address_6;
input 	onchip_memory2_0_s2_address_7;
input 	onchip_memory2_0_s2_address_8;
input 	onchip_memory2_0_s2_address_9;
input 	onchip_memory2_0_s2_address_10;
input 	onchip_memory2_0_s2_address_11;
input 	onchip_memory2_0_s2_address_12;
input 	onchip_memory2_0_s2_byteenable_0;
input 	onchip_memory2_0_s1_writedata_1;
input 	onchip_memory2_0_s2_writedata_1;
input 	onchip_memory2_0_s1_writedata_2;
input 	onchip_memory2_0_s2_writedata_2;
input 	onchip_memory2_0_s1_writedata_3;
input 	onchip_memory2_0_s2_writedata_3;
input 	onchip_memory2_0_s1_writedata_4;
input 	onchip_memory2_0_s2_writedata_4;
input 	onchip_memory2_0_s1_writedata_5;
input 	onchip_memory2_0_s2_writedata_5;
input 	onchip_memory2_0_s1_writedata_6;
input 	onchip_memory2_0_s2_writedata_6;
input 	onchip_memory2_0_s1_writedata_7;
input 	onchip_memory2_0_s2_writedata_7;
input 	onchip_memory2_0_s1_writedata_8;
input 	onchip_memory2_0_s1_byteenable_1;
input 	onchip_memory2_0_s2_writedata_8;
input 	onchip_memory2_0_s2_byteenable_1;
input 	onchip_memory2_0_s1_writedata_9;
input 	onchip_memory2_0_s2_writedata_9;
input 	onchip_memory2_0_s1_writedata_10;
input 	onchip_memory2_0_s2_writedata_10;
input 	onchip_memory2_0_s1_writedata_11;
input 	onchip_memory2_0_s2_writedata_11;
input 	onchip_memory2_0_s1_writedata_12;
input 	onchip_memory2_0_s2_writedata_12;
input 	onchip_memory2_0_s1_writedata_13;
input 	onchip_memory2_0_s2_writedata_13;
input 	onchip_memory2_0_s1_writedata_14;
input 	onchip_memory2_0_s2_writedata_14;
input 	onchip_memory2_0_s1_writedata_15;
input 	onchip_memory2_0_s2_writedata_15;
input 	onchip_memory2_0_s1_writedata_16;
input 	onchip_memory2_0_s1_byteenable_2;
input 	onchip_memory2_0_s2_writedata_16;
input 	onchip_memory2_0_s2_byteenable_2;
input 	onchip_memory2_0_s1_writedata_17;
input 	onchip_memory2_0_s2_writedata_17;
input 	onchip_memory2_0_s1_writedata_18;
input 	onchip_memory2_0_s2_writedata_18;
input 	onchip_memory2_0_s1_writedata_19;
input 	onchip_memory2_0_s2_writedata_19;
input 	onchip_memory2_0_s1_writedata_20;
input 	onchip_memory2_0_s2_writedata_20;
input 	onchip_memory2_0_s1_writedata_21;
input 	onchip_memory2_0_s2_writedata_21;
input 	onchip_memory2_0_s1_writedata_22;
input 	onchip_memory2_0_s2_writedata_22;
input 	onchip_memory2_0_s1_writedata_23;
input 	onchip_memory2_0_s2_writedata_23;
input 	onchip_memory2_0_s1_writedata_24;
input 	onchip_memory2_0_s1_byteenable_3;
input 	onchip_memory2_0_s2_writedata_24;
input 	onchip_memory2_0_s2_byteenable_3;
input 	onchip_memory2_0_s1_writedata_25;
input 	onchip_memory2_0_s2_writedata_25;
input 	onchip_memory2_0_s1_writedata_26;
input 	onchip_memory2_0_s2_writedata_26;
input 	onchip_memory2_0_s1_writedata_27;
input 	onchip_memory2_0_s2_writedata_27;
input 	onchip_memory2_0_s1_writedata_28;
input 	onchip_memory2_0_s2_writedata_28;
input 	onchip_memory2_0_s1_writedata_29;
input 	onchip_memory2_0_s2_writedata_29;
input 	onchip_memory2_0_s1_writedata_30;
input 	onchip_memory2_0_s2_writedata_30;
input 	onchip_memory2_0_s1_writedata_31;
input 	onchip_memory2_0_s2_writedata_31;
input 	onchip_memory2_0_s1_writedata_32;
input 	onchip_memory2_0_s1_byteenable_4;
input 	onchip_memory2_0_s2_writedata_32;
input 	onchip_memory2_0_s2_byteenable_4;
input 	onchip_memory2_0_s1_writedata_33;
input 	onchip_memory2_0_s2_writedata_33;
input 	onchip_memory2_0_s1_writedata_34;
input 	onchip_memory2_0_s2_writedata_34;
input 	onchip_memory2_0_s1_writedata_35;
input 	onchip_memory2_0_s2_writedata_35;
input 	onchip_memory2_0_s1_writedata_36;
input 	onchip_memory2_0_s2_writedata_36;
input 	onchip_memory2_0_s1_writedata_37;
input 	onchip_memory2_0_s2_writedata_37;
input 	onchip_memory2_0_s1_writedata_38;
input 	onchip_memory2_0_s2_writedata_38;
input 	onchip_memory2_0_s1_writedata_39;
input 	onchip_memory2_0_s2_writedata_39;
input 	onchip_memory2_0_s1_writedata_40;
input 	onchip_memory2_0_s1_byteenable_5;
input 	onchip_memory2_0_s2_writedata_40;
input 	onchip_memory2_0_s2_byteenable_5;
input 	onchip_memory2_0_s1_writedata_41;
input 	onchip_memory2_0_s2_writedata_41;
input 	onchip_memory2_0_s1_writedata_42;
input 	onchip_memory2_0_s2_writedata_42;
input 	onchip_memory2_0_s1_writedata_43;
input 	onchip_memory2_0_s2_writedata_43;
input 	onchip_memory2_0_s1_writedata_44;
input 	onchip_memory2_0_s2_writedata_44;
input 	onchip_memory2_0_s1_writedata_45;
input 	onchip_memory2_0_s2_writedata_45;
input 	onchip_memory2_0_s1_writedata_46;
input 	onchip_memory2_0_s2_writedata_46;
input 	onchip_memory2_0_s1_writedata_47;
input 	onchip_memory2_0_s2_writedata_47;
input 	onchip_memory2_0_s1_writedata_48;
input 	onchip_memory2_0_s1_byteenable_6;
input 	onchip_memory2_0_s2_writedata_48;
input 	onchip_memory2_0_s2_byteenable_6;
input 	onchip_memory2_0_s1_writedata_49;
input 	onchip_memory2_0_s2_writedata_49;
input 	onchip_memory2_0_s1_writedata_50;
input 	onchip_memory2_0_s2_writedata_50;
input 	onchip_memory2_0_s1_writedata_51;
input 	onchip_memory2_0_s2_writedata_51;
input 	onchip_memory2_0_s1_writedata_52;
input 	onchip_memory2_0_s2_writedata_52;
input 	onchip_memory2_0_s1_writedata_53;
input 	onchip_memory2_0_s2_writedata_53;
input 	onchip_memory2_0_s1_writedata_54;
input 	onchip_memory2_0_s2_writedata_54;
input 	onchip_memory2_0_s1_writedata_55;
input 	onchip_memory2_0_s2_writedata_55;
input 	onchip_memory2_0_s1_writedata_56;
input 	onchip_memory2_0_s1_byteenable_7;
input 	onchip_memory2_0_s2_writedata_56;
input 	onchip_memory2_0_s2_byteenable_7;
input 	onchip_memory2_0_s1_writedata_57;
input 	onchip_memory2_0_s2_writedata_57;
input 	onchip_memory2_0_s1_writedata_58;
input 	onchip_memory2_0_s2_writedata_58;
input 	onchip_memory2_0_s1_writedata_59;
input 	onchip_memory2_0_s2_writedata_59;
input 	onchip_memory2_0_s1_writedata_60;
input 	onchip_memory2_0_s2_writedata_60;
input 	onchip_memory2_0_s1_writedata_61;
input 	onchip_memory2_0_s2_writedata_61;
input 	onchip_memory2_0_s1_writedata_62;
input 	onchip_memory2_0_s2_writedata_62;
input 	onchip_memory2_0_s1_writedata_63;
input 	onchip_memory2_0_s2_writedata_63;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \clocken0~combout ;
wire \clocken1~combout ;


qtestpd_altsyncram_1 the_altsyncram(
	.result_node_0(result_node_0),
	.result_node_1(result_node_1),
	.result_node_2(result_node_2),
	.result_node_3(result_node_3),
	.result_node_4(result_node_4),
	.result_node_5(result_node_5),
	.result_node_6(result_node_6),
	.result_node_7(result_node_7),
	.result_node_8(result_node_8),
	.result_node_9(result_node_9),
	.result_node_10(result_node_10),
	.result_node_11(result_node_11),
	.result_node_12(result_node_12),
	.result_node_13(result_node_13),
	.result_node_14(result_node_14),
	.result_node_15(result_node_15),
	.result_node_16(result_node_16),
	.result_node_17(result_node_17),
	.result_node_18(result_node_18),
	.result_node_19(result_node_19),
	.result_node_20(result_node_20),
	.result_node_21(result_node_21),
	.result_node_22(result_node_22),
	.result_node_23(result_node_23),
	.result_node_24(result_node_24),
	.result_node_25(result_node_25),
	.result_node_26(result_node_26),
	.result_node_27(result_node_27),
	.result_node_28(result_node_28),
	.result_node_29(result_node_29),
	.result_node_30(result_node_30),
	.result_node_31(result_node_31),
	.result_node_32(result_node_32),
	.result_node_33(result_node_33),
	.result_node_34(result_node_34),
	.result_node_35(result_node_35),
	.result_node_36(result_node_36),
	.result_node_37(result_node_37),
	.result_node_38(result_node_38),
	.result_node_39(result_node_39),
	.result_node_40(result_node_40),
	.result_node_41(result_node_41),
	.result_node_42(result_node_42),
	.result_node_43(result_node_43),
	.result_node_44(result_node_44),
	.result_node_45(result_node_45),
	.result_node_46(result_node_46),
	.result_node_47(result_node_47),
	.result_node_48(result_node_48),
	.result_node_49(result_node_49),
	.result_node_50(result_node_50),
	.result_node_51(result_node_51),
	.result_node_52(result_node_52),
	.result_node_53(result_node_53),
	.result_node_54(result_node_54),
	.result_node_55(result_node_55),
	.result_node_56(result_node_56),
	.result_node_57(result_node_57),
	.result_node_58(result_node_58),
	.result_node_59(result_node_59),
	.result_node_60(result_node_60),
	.result_node_61(result_node_61),
	.result_node_62(result_node_62),
	.result_node_63(result_node_63),
	.result_node_01(result_node_01),
	.result_node_110(result_node_110),
	.result_node_210(result_node_210),
	.result_node_310(result_node_310),
	.result_node_410(result_node_410),
	.result_node_510(result_node_510),
	.result_node_64(result_node_64),
	.result_node_71(result_node_71),
	.result_node_81(result_node_81),
	.result_node_91(result_node_91),
	.result_node_101(result_node_101),
	.result_node_111(result_node_111),
	.result_node_121(result_node_121),
	.result_node_131(result_node_131),
	.result_node_141(result_node_141),
	.result_node_151(result_node_151),
	.result_node_161(result_node_161),
	.result_node_171(result_node_171),
	.result_node_181(result_node_181),
	.result_node_191(result_node_191),
	.result_node_201(result_node_201),
	.result_node_211(result_node_211),
	.result_node_221(result_node_221),
	.result_node_231(result_node_231),
	.result_node_241(result_node_241),
	.result_node_251(result_node_251),
	.result_node_261(result_node_261),
	.result_node_271(result_node_271),
	.result_node_281(result_node_281),
	.result_node_291(result_node_291),
	.result_node_301(result_node_301),
	.result_node_311(result_node_311),
	.result_node_321(result_node_321),
	.result_node_331(result_node_331),
	.result_node_341(result_node_341),
	.result_node_351(result_node_351),
	.result_node_361(result_node_361),
	.result_node_371(result_node_371),
	.result_node_381(result_node_381),
	.result_node_391(result_node_391),
	.result_node_401(result_node_401),
	.result_node_411(result_node_411),
	.result_node_421(result_node_421),
	.result_node_431(result_node_431),
	.result_node_441(result_node_441),
	.result_node_451(result_node_451),
	.result_node_461(result_node_461),
	.result_node_471(result_node_471),
	.result_node_481(result_node_481),
	.result_node_491(result_node_491),
	.result_node_501(result_node_501),
	.result_node_511(result_node_511),
	.result_node_521(result_node_521),
	.result_node_531(result_node_531),
	.result_node_541(result_node_541),
	.result_node_551(result_node_551),
	.result_node_561(result_node_561),
	.result_node_571(result_node_571),
	.result_node_581(result_node_581),
	.result_node_591(result_node_591),
	.result_node_601(result_node_601),
	.result_node_611(result_node_611),
	.result_node_621(result_node_621),
	.result_node_631(result_node_631),
	.clocken0(\clocken0~combout ),
	.clocken1(\clocken1~combout ),
	.address_a({onchip_memory2_0_s1_address_13,onchip_memory2_0_s1_address_12,onchip_memory2_0_s1_address_11,onchip_memory2_0_s1_address_10,onchip_memory2_0_s1_address_9,onchip_memory2_0_s1_address_8,onchip_memory2_0_s1_address_7,onchip_memory2_0_s1_address_6,
onchip_memory2_0_s1_address_5,onchip_memory2_0_s1_address_4,onchip_memory2_0_s1_address_3,onchip_memory2_0_s1_address_2,onchip_memory2_0_s1_address_1,onchip_memory2_0_s1_address_0}),
	.onchip_memory2_0_s1_chipselect(onchip_memory2_0_s1_chipselect),
	.onchip_memory2_0_s1_write(onchip_memory2_0_s1_write),
	.address_b({onchip_memory2_0_s2_address_13,onchip_memory2_0_s2_address_12,onchip_memory2_0_s2_address_11,onchip_memory2_0_s2_address_10,onchip_memory2_0_s2_address_9,onchip_memory2_0_s2_address_8,onchip_memory2_0_s2_address_7,onchip_memory2_0_s2_address_6,
onchip_memory2_0_s2_address_5,onchip_memory2_0_s2_address_4,onchip_memory2_0_s2_address_3,onchip_memory2_0_s2_address_2,onchip_memory2_0_s2_address_1,onchip_memory2_0_s2_address_0}),
	.onchip_memory2_0_s2_chipselect(onchip_memory2_0_s2_chipselect),
	.onchip_memory2_0_s2_write(onchip_memory2_0_s2_write),
	.clock1(clk_clk),
	.data_a({onchip_memory2_0_s1_writedata_63,onchip_memory2_0_s1_writedata_62,onchip_memory2_0_s1_writedata_61,onchip_memory2_0_s1_writedata_60,onchip_memory2_0_s1_writedata_59,onchip_memory2_0_s1_writedata_58,onchip_memory2_0_s1_writedata_57,onchip_memory2_0_s1_writedata_56,
onchip_memory2_0_s1_writedata_55,onchip_memory2_0_s1_writedata_54,onchip_memory2_0_s1_writedata_53,onchip_memory2_0_s1_writedata_52,onchip_memory2_0_s1_writedata_51,onchip_memory2_0_s1_writedata_50,onchip_memory2_0_s1_writedata_49,onchip_memory2_0_s1_writedata_48,
onchip_memory2_0_s1_writedata_47,onchip_memory2_0_s1_writedata_46,onchip_memory2_0_s1_writedata_45,onchip_memory2_0_s1_writedata_44,onchip_memory2_0_s1_writedata_43,onchip_memory2_0_s1_writedata_42,onchip_memory2_0_s1_writedata_41,onchip_memory2_0_s1_writedata_40,
onchip_memory2_0_s1_writedata_39,onchip_memory2_0_s1_writedata_38,onchip_memory2_0_s1_writedata_37,onchip_memory2_0_s1_writedata_36,onchip_memory2_0_s1_writedata_35,onchip_memory2_0_s1_writedata_34,onchip_memory2_0_s1_writedata_33,onchip_memory2_0_s1_writedata_32,
onchip_memory2_0_s1_writedata_31,onchip_memory2_0_s1_writedata_30,onchip_memory2_0_s1_writedata_29,onchip_memory2_0_s1_writedata_28,onchip_memory2_0_s1_writedata_27,onchip_memory2_0_s1_writedata_26,onchip_memory2_0_s1_writedata_25,onchip_memory2_0_s1_writedata_24,
onchip_memory2_0_s1_writedata_23,onchip_memory2_0_s1_writedata_22,onchip_memory2_0_s1_writedata_21,onchip_memory2_0_s1_writedata_20,onchip_memory2_0_s1_writedata_19,onchip_memory2_0_s1_writedata_18,onchip_memory2_0_s1_writedata_17,onchip_memory2_0_s1_writedata_16,
onchip_memory2_0_s1_writedata_15,onchip_memory2_0_s1_writedata_14,onchip_memory2_0_s1_writedata_13,onchip_memory2_0_s1_writedata_12,onchip_memory2_0_s1_writedata_11,onchip_memory2_0_s1_writedata_10,onchip_memory2_0_s1_writedata_9,onchip_memory2_0_s1_writedata_8,
onchip_memory2_0_s1_writedata_7,onchip_memory2_0_s1_writedata_6,onchip_memory2_0_s1_writedata_5,onchip_memory2_0_s1_writedata_4,onchip_memory2_0_s1_writedata_3,onchip_memory2_0_s1_writedata_2,onchip_memory2_0_s1_writedata_1,onchip_memory2_0_s1_writedata_0}),
	.byteena_a({onchip_memory2_0_s1_byteenable_7,onchip_memory2_0_s1_byteenable_6,onchip_memory2_0_s1_byteenable_5,onchip_memory2_0_s1_byteenable_4,onchip_memory2_0_s1_byteenable_3,onchip_memory2_0_s1_byteenable_2,onchip_memory2_0_s1_byteenable_1,onchip_memory2_0_s1_byteenable_0}),
	.data_b({onchip_memory2_0_s2_writedata_63,onchip_memory2_0_s2_writedata_62,onchip_memory2_0_s2_writedata_61,onchip_memory2_0_s2_writedata_60,onchip_memory2_0_s2_writedata_59,onchip_memory2_0_s2_writedata_58,onchip_memory2_0_s2_writedata_57,onchip_memory2_0_s2_writedata_56,
onchip_memory2_0_s2_writedata_55,onchip_memory2_0_s2_writedata_54,onchip_memory2_0_s2_writedata_53,onchip_memory2_0_s2_writedata_52,onchip_memory2_0_s2_writedata_51,onchip_memory2_0_s2_writedata_50,onchip_memory2_0_s2_writedata_49,onchip_memory2_0_s2_writedata_48,
onchip_memory2_0_s2_writedata_47,onchip_memory2_0_s2_writedata_46,onchip_memory2_0_s2_writedata_45,onchip_memory2_0_s2_writedata_44,onchip_memory2_0_s2_writedata_43,onchip_memory2_0_s2_writedata_42,onchip_memory2_0_s2_writedata_41,onchip_memory2_0_s2_writedata_40,
onchip_memory2_0_s2_writedata_39,onchip_memory2_0_s2_writedata_38,onchip_memory2_0_s2_writedata_37,onchip_memory2_0_s2_writedata_36,onchip_memory2_0_s2_writedata_35,onchip_memory2_0_s2_writedata_34,onchip_memory2_0_s2_writedata_33,onchip_memory2_0_s2_writedata_32,
onchip_memory2_0_s2_writedata_31,onchip_memory2_0_s2_writedata_30,onchip_memory2_0_s2_writedata_29,onchip_memory2_0_s2_writedata_28,onchip_memory2_0_s2_writedata_27,onchip_memory2_0_s2_writedata_26,onchip_memory2_0_s2_writedata_25,onchip_memory2_0_s2_writedata_24,
onchip_memory2_0_s2_writedata_23,onchip_memory2_0_s2_writedata_22,onchip_memory2_0_s2_writedata_21,onchip_memory2_0_s2_writedata_20,onchip_memory2_0_s2_writedata_19,onchip_memory2_0_s2_writedata_18,onchip_memory2_0_s2_writedata_17,onchip_memory2_0_s2_writedata_16,
onchip_memory2_0_s2_writedata_15,onchip_memory2_0_s2_writedata_14,onchip_memory2_0_s2_writedata_13,onchip_memory2_0_s2_writedata_12,onchip_memory2_0_s2_writedata_11,onchip_memory2_0_s2_writedata_10,onchip_memory2_0_s2_writedata_9,onchip_memory2_0_s2_writedata_8,
onchip_memory2_0_s2_writedata_7,onchip_memory2_0_s2_writedata_6,onchip_memory2_0_s2_writedata_5,onchip_memory2_0_s2_writedata_4,onchip_memory2_0_s2_writedata_3,onchip_memory2_0_s2_writedata_2,onchip_memory2_0_s2_writedata_1,onchip_memory2_0_s2_writedata_0}),
	.byteena_b({onchip_memory2_0_s2_byteenable_7,onchip_memory2_0_s2_byteenable_6,onchip_memory2_0_s2_byteenable_5,onchip_memory2_0_s2_byteenable_4,onchip_memory2_0_s2_byteenable_3,onchip_memory2_0_s2_byteenable_2,onchip_memory2_0_s2_byteenable_1,onchip_memory2_0_s2_byteenable_0}));

cycloneiv_lcell_comb clocken0(
	.dataa(onchip_memory2_0_s1_clken),
	.datab(gnd),
	.datac(gnd),
	.datad(r_early_rst),
	.cin(gnd),
	.combout(\clocken0~combout ),
	.cout());
defparam clocken0.lut_mask = 16'h00AA;
defparam clocken0.sum_lutc_input = "datac";

cycloneiv_lcell_comb clocken1(
	.dataa(onchip_memory2_0_s2_clken),
	.datab(gnd),
	.datac(gnd),
	.datad(r_early_rst),
	.cin(gnd),
	.combout(\clocken1~combout ),
	.cout());
defparam clocken1.lut_mask = 16'h00AA;
defparam clocken1.sum_lutc_input = "datac";

endmodule

module qtestpd_altsyncram_1 (
	result_node_0,
	result_node_1,
	result_node_2,
	result_node_3,
	result_node_4,
	result_node_5,
	result_node_6,
	result_node_7,
	result_node_8,
	result_node_9,
	result_node_10,
	result_node_11,
	result_node_12,
	result_node_13,
	result_node_14,
	result_node_15,
	result_node_16,
	result_node_17,
	result_node_18,
	result_node_19,
	result_node_20,
	result_node_21,
	result_node_22,
	result_node_23,
	result_node_24,
	result_node_25,
	result_node_26,
	result_node_27,
	result_node_28,
	result_node_29,
	result_node_30,
	result_node_31,
	result_node_32,
	result_node_33,
	result_node_34,
	result_node_35,
	result_node_36,
	result_node_37,
	result_node_38,
	result_node_39,
	result_node_40,
	result_node_41,
	result_node_42,
	result_node_43,
	result_node_44,
	result_node_45,
	result_node_46,
	result_node_47,
	result_node_48,
	result_node_49,
	result_node_50,
	result_node_51,
	result_node_52,
	result_node_53,
	result_node_54,
	result_node_55,
	result_node_56,
	result_node_57,
	result_node_58,
	result_node_59,
	result_node_60,
	result_node_61,
	result_node_62,
	result_node_63,
	result_node_01,
	result_node_110,
	result_node_210,
	result_node_310,
	result_node_410,
	result_node_510,
	result_node_64,
	result_node_71,
	result_node_81,
	result_node_91,
	result_node_101,
	result_node_111,
	result_node_121,
	result_node_131,
	result_node_141,
	result_node_151,
	result_node_161,
	result_node_171,
	result_node_181,
	result_node_191,
	result_node_201,
	result_node_211,
	result_node_221,
	result_node_231,
	result_node_241,
	result_node_251,
	result_node_261,
	result_node_271,
	result_node_281,
	result_node_291,
	result_node_301,
	result_node_311,
	result_node_321,
	result_node_331,
	result_node_341,
	result_node_351,
	result_node_361,
	result_node_371,
	result_node_381,
	result_node_391,
	result_node_401,
	result_node_411,
	result_node_421,
	result_node_431,
	result_node_441,
	result_node_451,
	result_node_461,
	result_node_471,
	result_node_481,
	result_node_491,
	result_node_501,
	result_node_511,
	result_node_521,
	result_node_531,
	result_node_541,
	result_node_551,
	result_node_561,
	result_node_571,
	result_node_581,
	result_node_591,
	result_node_601,
	result_node_611,
	result_node_621,
	result_node_631,
	clocken0,
	clocken1,
	address_a,
	onchip_memory2_0_s1_chipselect,
	onchip_memory2_0_s1_write,
	address_b,
	onchip_memory2_0_s2_chipselect,
	onchip_memory2_0_s2_write,
	clock1,
	data_a,
	byteena_a,
	data_b,
	byteena_b)/* synthesis synthesis_greybox=0 */;
output 	result_node_0;
output 	result_node_1;
output 	result_node_2;
output 	result_node_3;
output 	result_node_4;
output 	result_node_5;
output 	result_node_6;
output 	result_node_7;
output 	result_node_8;
output 	result_node_9;
output 	result_node_10;
output 	result_node_11;
output 	result_node_12;
output 	result_node_13;
output 	result_node_14;
output 	result_node_15;
output 	result_node_16;
output 	result_node_17;
output 	result_node_18;
output 	result_node_19;
output 	result_node_20;
output 	result_node_21;
output 	result_node_22;
output 	result_node_23;
output 	result_node_24;
output 	result_node_25;
output 	result_node_26;
output 	result_node_27;
output 	result_node_28;
output 	result_node_29;
output 	result_node_30;
output 	result_node_31;
output 	result_node_32;
output 	result_node_33;
output 	result_node_34;
output 	result_node_35;
output 	result_node_36;
output 	result_node_37;
output 	result_node_38;
output 	result_node_39;
output 	result_node_40;
output 	result_node_41;
output 	result_node_42;
output 	result_node_43;
output 	result_node_44;
output 	result_node_45;
output 	result_node_46;
output 	result_node_47;
output 	result_node_48;
output 	result_node_49;
output 	result_node_50;
output 	result_node_51;
output 	result_node_52;
output 	result_node_53;
output 	result_node_54;
output 	result_node_55;
output 	result_node_56;
output 	result_node_57;
output 	result_node_58;
output 	result_node_59;
output 	result_node_60;
output 	result_node_61;
output 	result_node_62;
output 	result_node_63;
output 	result_node_01;
output 	result_node_110;
output 	result_node_210;
output 	result_node_310;
output 	result_node_410;
output 	result_node_510;
output 	result_node_64;
output 	result_node_71;
output 	result_node_81;
output 	result_node_91;
output 	result_node_101;
output 	result_node_111;
output 	result_node_121;
output 	result_node_131;
output 	result_node_141;
output 	result_node_151;
output 	result_node_161;
output 	result_node_171;
output 	result_node_181;
output 	result_node_191;
output 	result_node_201;
output 	result_node_211;
output 	result_node_221;
output 	result_node_231;
output 	result_node_241;
output 	result_node_251;
output 	result_node_261;
output 	result_node_271;
output 	result_node_281;
output 	result_node_291;
output 	result_node_301;
output 	result_node_311;
output 	result_node_321;
output 	result_node_331;
output 	result_node_341;
output 	result_node_351;
output 	result_node_361;
output 	result_node_371;
output 	result_node_381;
output 	result_node_391;
output 	result_node_401;
output 	result_node_411;
output 	result_node_421;
output 	result_node_431;
output 	result_node_441;
output 	result_node_451;
output 	result_node_461;
output 	result_node_471;
output 	result_node_481;
output 	result_node_491;
output 	result_node_501;
output 	result_node_511;
output 	result_node_521;
output 	result_node_531;
output 	result_node_541;
output 	result_node_551;
output 	result_node_561;
output 	result_node_571;
output 	result_node_581;
output 	result_node_591;
output 	result_node_601;
output 	result_node_611;
output 	result_node_621;
output 	result_node_631;
input 	clocken0;
input 	clocken1;
input 	[13:0] address_a;
input 	onchip_memory2_0_s1_chipselect;
input 	onchip_memory2_0_s1_write;
input 	[13:0] address_b;
input 	onchip_memory2_0_s2_chipselect;
input 	onchip_memory2_0_s2_write;
input 	clock1;
input 	[63:0] data_a;
input 	[7:0] byteena_a;
input 	[63:0] data_b;
input 	[7:0] byteena_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



qtestpd_altsyncram_6342 auto_generated(
	.result_node_0(result_node_0),
	.result_node_1(result_node_1),
	.result_node_2(result_node_2),
	.result_node_3(result_node_3),
	.result_node_4(result_node_4),
	.result_node_5(result_node_5),
	.result_node_6(result_node_6),
	.result_node_7(result_node_7),
	.result_node_8(result_node_8),
	.result_node_9(result_node_9),
	.result_node_10(result_node_10),
	.result_node_11(result_node_11),
	.result_node_12(result_node_12),
	.result_node_13(result_node_13),
	.result_node_14(result_node_14),
	.result_node_15(result_node_15),
	.result_node_16(result_node_16),
	.result_node_17(result_node_17),
	.result_node_18(result_node_18),
	.result_node_19(result_node_19),
	.result_node_20(result_node_20),
	.result_node_21(result_node_21),
	.result_node_22(result_node_22),
	.result_node_23(result_node_23),
	.result_node_24(result_node_24),
	.result_node_25(result_node_25),
	.result_node_26(result_node_26),
	.result_node_27(result_node_27),
	.result_node_28(result_node_28),
	.result_node_29(result_node_29),
	.result_node_30(result_node_30),
	.result_node_31(result_node_31),
	.result_node_32(result_node_32),
	.result_node_33(result_node_33),
	.result_node_34(result_node_34),
	.result_node_35(result_node_35),
	.result_node_36(result_node_36),
	.result_node_37(result_node_37),
	.result_node_38(result_node_38),
	.result_node_39(result_node_39),
	.result_node_40(result_node_40),
	.result_node_41(result_node_41),
	.result_node_42(result_node_42),
	.result_node_43(result_node_43),
	.result_node_44(result_node_44),
	.result_node_45(result_node_45),
	.result_node_46(result_node_46),
	.result_node_47(result_node_47),
	.result_node_48(result_node_48),
	.result_node_49(result_node_49),
	.result_node_50(result_node_50),
	.result_node_51(result_node_51),
	.result_node_52(result_node_52),
	.result_node_53(result_node_53),
	.result_node_54(result_node_54),
	.result_node_55(result_node_55),
	.result_node_56(result_node_56),
	.result_node_57(result_node_57),
	.result_node_58(result_node_58),
	.result_node_59(result_node_59),
	.result_node_60(result_node_60),
	.result_node_61(result_node_61),
	.result_node_62(result_node_62),
	.result_node_63(result_node_63),
	.result_node_01(result_node_01),
	.result_node_110(result_node_110),
	.result_node_210(result_node_210),
	.result_node_310(result_node_310),
	.result_node_410(result_node_410),
	.result_node_510(result_node_510),
	.result_node_64(result_node_64),
	.result_node_71(result_node_71),
	.result_node_81(result_node_81),
	.result_node_91(result_node_91),
	.result_node_101(result_node_101),
	.result_node_111(result_node_111),
	.result_node_121(result_node_121),
	.result_node_131(result_node_131),
	.result_node_141(result_node_141),
	.result_node_151(result_node_151),
	.result_node_161(result_node_161),
	.result_node_171(result_node_171),
	.result_node_181(result_node_181),
	.result_node_191(result_node_191),
	.result_node_201(result_node_201),
	.result_node_211(result_node_211),
	.result_node_221(result_node_221),
	.result_node_231(result_node_231),
	.result_node_241(result_node_241),
	.result_node_251(result_node_251),
	.result_node_261(result_node_261),
	.result_node_271(result_node_271),
	.result_node_281(result_node_281),
	.result_node_291(result_node_291),
	.result_node_301(result_node_301),
	.result_node_311(result_node_311),
	.result_node_321(result_node_321),
	.result_node_331(result_node_331),
	.result_node_341(result_node_341),
	.result_node_351(result_node_351),
	.result_node_361(result_node_361),
	.result_node_371(result_node_371),
	.result_node_381(result_node_381),
	.result_node_391(result_node_391),
	.result_node_401(result_node_401),
	.result_node_411(result_node_411),
	.result_node_421(result_node_421),
	.result_node_431(result_node_431),
	.result_node_441(result_node_441),
	.result_node_451(result_node_451),
	.result_node_461(result_node_461),
	.result_node_471(result_node_471),
	.result_node_481(result_node_481),
	.result_node_491(result_node_491),
	.result_node_501(result_node_501),
	.result_node_511(result_node_511),
	.result_node_521(result_node_521),
	.result_node_531(result_node_531),
	.result_node_541(result_node_541),
	.result_node_551(result_node_551),
	.result_node_561(result_node_561),
	.result_node_571(result_node_571),
	.result_node_581(result_node_581),
	.result_node_591(result_node_591),
	.result_node_601(result_node_601),
	.result_node_611(result_node_611),
	.result_node_621(result_node_621),
	.result_node_631(result_node_631),
	.clocken0(clocken0),
	.clocken1(clocken1),
	.address_a({address_a[13],address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.onchip_memory2_0_s1_chipselect(onchip_memory2_0_s1_chipselect),
	.onchip_memory2_0_s1_write(onchip_memory2_0_s1_write),
	.address_b({address_b[13],address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.onchip_memory2_0_s2_chipselect(onchip_memory2_0_s2_chipselect),
	.onchip_memory2_0_s2_write(onchip_memory2_0_s2_write),
	.clock1(clock1),
	.clock0(clock1),
	.data_a({data_a[63],data_a[62],data_a[61],data_a[60],data_a[59],data_a[58],data_a[57],data_a[56],data_a[55],data_a[54],data_a[53],data_a[52],data_a[51],data_a[50],data_a[49],data_a[48],data_a[47],data_a[46],data_a[45],data_a[44],data_a[43],data_a[42],data_a[41],data_a[40],data_a[39],data_a[38],data_a[37],data_a[36],data_a[35],data_a[34],data_a[33],data_a[32],data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],
data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.byteena_a({byteena_a[7],byteena_a[6],byteena_a[5],byteena_a[4],byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.data_b({data_b[63],data_b[62],data_b[61],data_b[60],data_b[59],data_b[58],data_b[57],data_b[56],data_b[55],data_b[54],data_b[53],data_b[52],data_b[51],data_b[50],data_b[49],data_b[48],data_b[47],data_b[46],data_b[45],data_b[44],data_b[43],data_b[42],data_b[41],data_b[40],data_b[39],data_b[38],data_b[37],data_b[36],data_b[35],data_b[34],data_b[33],data_b[32],data_b[31],data_b[30],data_b[29],data_b[28],data_b[27],data_b[26],data_b[25],data_b[24],data_b[23],data_b[22],
data_b[21],data_b[20],data_b[19],data_b[18],data_b[17],data_b[16],data_b[15],data_b[14],data_b[13],data_b[12],data_b[11],data_b[10],data_b[9],data_b[8],data_b[7],data_b[6],data_b[5],data_b[4],data_b[3],data_b[2],data_b[1],data_b[0]}),
	.byteena_b({byteena_b[7],byteena_b[6],byteena_b[5],byteena_b[4],byteena_b[3],byteena_b[2],byteena_b[1],byteena_b[0]}));

endmodule

module qtestpd_altsyncram_6342 (
	result_node_0,
	result_node_1,
	result_node_2,
	result_node_3,
	result_node_4,
	result_node_5,
	result_node_6,
	result_node_7,
	result_node_8,
	result_node_9,
	result_node_10,
	result_node_11,
	result_node_12,
	result_node_13,
	result_node_14,
	result_node_15,
	result_node_16,
	result_node_17,
	result_node_18,
	result_node_19,
	result_node_20,
	result_node_21,
	result_node_22,
	result_node_23,
	result_node_24,
	result_node_25,
	result_node_26,
	result_node_27,
	result_node_28,
	result_node_29,
	result_node_30,
	result_node_31,
	result_node_32,
	result_node_33,
	result_node_34,
	result_node_35,
	result_node_36,
	result_node_37,
	result_node_38,
	result_node_39,
	result_node_40,
	result_node_41,
	result_node_42,
	result_node_43,
	result_node_44,
	result_node_45,
	result_node_46,
	result_node_47,
	result_node_48,
	result_node_49,
	result_node_50,
	result_node_51,
	result_node_52,
	result_node_53,
	result_node_54,
	result_node_55,
	result_node_56,
	result_node_57,
	result_node_58,
	result_node_59,
	result_node_60,
	result_node_61,
	result_node_62,
	result_node_63,
	result_node_01,
	result_node_110,
	result_node_210,
	result_node_310,
	result_node_410,
	result_node_510,
	result_node_64,
	result_node_71,
	result_node_81,
	result_node_91,
	result_node_101,
	result_node_111,
	result_node_121,
	result_node_131,
	result_node_141,
	result_node_151,
	result_node_161,
	result_node_171,
	result_node_181,
	result_node_191,
	result_node_201,
	result_node_211,
	result_node_221,
	result_node_231,
	result_node_241,
	result_node_251,
	result_node_261,
	result_node_271,
	result_node_281,
	result_node_291,
	result_node_301,
	result_node_311,
	result_node_321,
	result_node_331,
	result_node_341,
	result_node_351,
	result_node_361,
	result_node_371,
	result_node_381,
	result_node_391,
	result_node_401,
	result_node_411,
	result_node_421,
	result_node_431,
	result_node_441,
	result_node_451,
	result_node_461,
	result_node_471,
	result_node_481,
	result_node_491,
	result_node_501,
	result_node_511,
	result_node_521,
	result_node_531,
	result_node_541,
	result_node_551,
	result_node_561,
	result_node_571,
	result_node_581,
	result_node_591,
	result_node_601,
	result_node_611,
	result_node_621,
	result_node_631,
	clocken0,
	clocken1,
	address_a,
	onchip_memory2_0_s1_chipselect,
	onchip_memory2_0_s1_write,
	address_b,
	onchip_memory2_0_s2_chipselect,
	onchip_memory2_0_s2_write,
	clock1,
	clock0,
	data_a,
	byteena_a,
	data_b,
	byteena_b)/* synthesis synthesis_greybox=0 */;
output 	result_node_0;
output 	result_node_1;
output 	result_node_2;
output 	result_node_3;
output 	result_node_4;
output 	result_node_5;
output 	result_node_6;
output 	result_node_7;
output 	result_node_8;
output 	result_node_9;
output 	result_node_10;
output 	result_node_11;
output 	result_node_12;
output 	result_node_13;
output 	result_node_14;
output 	result_node_15;
output 	result_node_16;
output 	result_node_17;
output 	result_node_18;
output 	result_node_19;
output 	result_node_20;
output 	result_node_21;
output 	result_node_22;
output 	result_node_23;
output 	result_node_24;
output 	result_node_25;
output 	result_node_26;
output 	result_node_27;
output 	result_node_28;
output 	result_node_29;
output 	result_node_30;
output 	result_node_31;
output 	result_node_32;
output 	result_node_33;
output 	result_node_34;
output 	result_node_35;
output 	result_node_36;
output 	result_node_37;
output 	result_node_38;
output 	result_node_39;
output 	result_node_40;
output 	result_node_41;
output 	result_node_42;
output 	result_node_43;
output 	result_node_44;
output 	result_node_45;
output 	result_node_46;
output 	result_node_47;
output 	result_node_48;
output 	result_node_49;
output 	result_node_50;
output 	result_node_51;
output 	result_node_52;
output 	result_node_53;
output 	result_node_54;
output 	result_node_55;
output 	result_node_56;
output 	result_node_57;
output 	result_node_58;
output 	result_node_59;
output 	result_node_60;
output 	result_node_61;
output 	result_node_62;
output 	result_node_63;
output 	result_node_01;
output 	result_node_110;
output 	result_node_210;
output 	result_node_310;
output 	result_node_410;
output 	result_node_510;
output 	result_node_64;
output 	result_node_71;
output 	result_node_81;
output 	result_node_91;
output 	result_node_101;
output 	result_node_111;
output 	result_node_121;
output 	result_node_131;
output 	result_node_141;
output 	result_node_151;
output 	result_node_161;
output 	result_node_171;
output 	result_node_181;
output 	result_node_191;
output 	result_node_201;
output 	result_node_211;
output 	result_node_221;
output 	result_node_231;
output 	result_node_241;
output 	result_node_251;
output 	result_node_261;
output 	result_node_271;
output 	result_node_281;
output 	result_node_291;
output 	result_node_301;
output 	result_node_311;
output 	result_node_321;
output 	result_node_331;
output 	result_node_341;
output 	result_node_351;
output 	result_node_361;
output 	result_node_371;
output 	result_node_381;
output 	result_node_391;
output 	result_node_401;
output 	result_node_411;
output 	result_node_421;
output 	result_node_431;
output 	result_node_441;
output 	result_node_451;
output 	result_node_461;
output 	result_node_471;
output 	result_node_481;
output 	result_node_491;
output 	result_node_501;
output 	result_node_511;
output 	result_node_521;
output 	result_node_531;
output 	result_node_541;
output 	result_node_551;
output 	result_node_561;
output 	result_node_571;
output 	result_node_581;
output 	result_node_591;
output 	result_node_601;
output 	result_node_611;
output 	result_node_621;
output 	result_node_631;
input 	clocken0;
input 	clocken1;
input 	[13:0] address_a;
input 	onchip_memory2_0_s1_chipselect;
input 	onchip_memory2_0_s1_write;
input 	[13:0] address_b;
input 	onchip_memory2_0_s2_chipselect;
input 	onchip_memory2_0_s2_write;
input 	clock1;
input 	clock0;
input 	[63:0] data_a;
input 	[7:0] byteena_a;
input 	[63:0] data_b;
input 	[7:0] byteena_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ram_block1a64~portadataout ;
wire \ram_block1a64~PORTBDATAOUT0 ;
wire \ram_block1a0~portadataout ;
wire \ram_block1a0~PORTBDATAOUT0 ;
wire \ram_block1a65~portadataout ;
wire \ram_block1a65~PORTBDATAOUT0 ;
wire \ram_block1a1~portadataout ;
wire \ram_block1a1~PORTBDATAOUT0 ;
wire \ram_block1a66~portadataout ;
wire \ram_block1a66~PORTBDATAOUT0 ;
wire \ram_block1a2~portadataout ;
wire \ram_block1a2~PORTBDATAOUT0 ;
wire \ram_block1a67~portadataout ;
wire \ram_block1a67~PORTBDATAOUT0 ;
wire \ram_block1a3~portadataout ;
wire \ram_block1a3~PORTBDATAOUT0 ;
wire \ram_block1a68~portadataout ;
wire \ram_block1a68~PORTBDATAOUT0 ;
wire \ram_block1a4~portadataout ;
wire \ram_block1a4~PORTBDATAOUT0 ;
wire \ram_block1a69~portadataout ;
wire \ram_block1a69~PORTBDATAOUT0 ;
wire \ram_block1a5~portadataout ;
wire \ram_block1a5~PORTBDATAOUT0 ;
wire \ram_block1a70~portadataout ;
wire \ram_block1a70~PORTBDATAOUT0 ;
wire \ram_block1a6~portadataout ;
wire \ram_block1a6~PORTBDATAOUT0 ;
wire \ram_block1a71~portadataout ;
wire \ram_block1a71~PORTBDATAOUT0 ;
wire \ram_block1a7~portadataout ;
wire \ram_block1a7~PORTBDATAOUT0 ;
wire \ram_block1a72~portadataout ;
wire \ram_block1a72~PORTBDATAOUT0 ;
wire \ram_block1a8~portadataout ;
wire \ram_block1a8~PORTBDATAOUT0 ;
wire \ram_block1a73~portadataout ;
wire \ram_block1a73~PORTBDATAOUT0 ;
wire \ram_block1a9~portadataout ;
wire \ram_block1a9~PORTBDATAOUT0 ;
wire \ram_block1a74~portadataout ;
wire \ram_block1a74~PORTBDATAOUT0 ;
wire \ram_block1a10~portadataout ;
wire \ram_block1a10~PORTBDATAOUT0 ;
wire \ram_block1a75~portadataout ;
wire \ram_block1a75~PORTBDATAOUT0 ;
wire \ram_block1a11~portadataout ;
wire \ram_block1a11~PORTBDATAOUT0 ;
wire \ram_block1a76~portadataout ;
wire \ram_block1a76~PORTBDATAOUT0 ;
wire \ram_block1a12~portadataout ;
wire \ram_block1a12~PORTBDATAOUT0 ;
wire \ram_block1a77~portadataout ;
wire \ram_block1a77~PORTBDATAOUT0 ;
wire \ram_block1a13~portadataout ;
wire \ram_block1a13~PORTBDATAOUT0 ;
wire \ram_block1a78~portadataout ;
wire \ram_block1a78~PORTBDATAOUT0 ;
wire \ram_block1a14~portadataout ;
wire \ram_block1a14~PORTBDATAOUT0 ;
wire \ram_block1a79~portadataout ;
wire \ram_block1a79~PORTBDATAOUT0 ;
wire \ram_block1a15~portadataout ;
wire \ram_block1a15~PORTBDATAOUT0 ;
wire \ram_block1a80~portadataout ;
wire \ram_block1a80~PORTBDATAOUT0 ;
wire \ram_block1a16~portadataout ;
wire \ram_block1a16~PORTBDATAOUT0 ;
wire \ram_block1a81~portadataout ;
wire \ram_block1a81~PORTBDATAOUT0 ;
wire \ram_block1a17~portadataout ;
wire \ram_block1a17~PORTBDATAOUT0 ;
wire \ram_block1a82~portadataout ;
wire \ram_block1a82~PORTBDATAOUT0 ;
wire \ram_block1a18~portadataout ;
wire \ram_block1a18~PORTBDATAOUT0 ;
wire \ram_block1a83~portadataout ;
wire \ram_block1a83~PORTBDATAOUT0 ;
wire \ram_block1a19~portadataout ;
wire \ram_block1a19~PORTBDATAOUT0 ;
wire \ram_block1a84~portadataout ;
wire \ram_block1a84~PORTBDATAOUT0 ;
wire \ram_block1a20~portadataout ;
wire \ram_block1a20~PORTBDATAOUT0 ;
wire \ram_block1a85~portadataout ;
wire \ram_block1a85~PORTBDATAOUT0 ;
wire \ram_block1a21~portadataout ;
wire \ram_block1a21~PORTBDATAOUT0 ;
wire \ram_block1a86~portadataout ;
wire \ram_block1a86~PORTBDATAOUT0 ;
wire \ram_block1a22~portadataout ;
wire \ram_block1a22~PORTBDATAOUT0 ;
wire \ram_block1a87~portadataout ;
wire \ram_block1a87~PORTBDATAOUT0 ;
wire \ram_block1a23~portadataout ;
wire \ram_block1a23~PORTBDATAOUT0 ;
wire \ram_block1a88~portadataout ;
wire \ram_block1a88~PORTBDATAOUT0 ;
wire \ram_block1a24~portadataout ;
wire \ram_block1a24~PORTBDATAOUT0 ;
wire \ram_block1a89~portadataout ;
wire \ram_block1a89~PORTBDATAOUT0 ;
wire \ram_block1a25~portadataout ;
wire \ram_block1a25~PORTBDATAOUT0 ;
wire \ram_block1a90~portadataout ;
wire \ram_block1a90~PORTBDATAOUT0 ;
wire \ram_block1a26~portadataout ;
wire \ram_block1a26~PORTBDATAOUT0 ;
wire \ram_block1a91~portadataout ;
wire \ram_block1a91~PORTBDATAOUT0 ;
wire \ram_block1a27~portadataout ;
wire \ram_block1a27~PORTBDATAOUT0 ;
wire \ram_block1a92~portadataout ;
wire \ram_block1a92~PORTBDATAOUT0 ;
wire \ram_block1a28~portadataout ;
wire \ram_block1a28~PORTBDATAOUT0 ;
wire \ram_block1a93~portadataout ;
wire \ram_block1a93~PORTBDATAOUT0 ;
wire \ram_block1a29~portadataout ;
wire \ram_block1a29~PORTBDATAOUT0 ;
wire \ram_block1a94~portadataout ;
wire \ram_block1a94~PORTBDATAOUT0 ;
wire \ram_block1a30~portadataout ;
wire \ram_block1a30~PORTBDATAOUT0 ;
wire \ram_block1a95~portadataout ;
wire \ram_block1a95~PORTBDATAOUT0 ;
wire \ram_block1a31~portadataout ;
wire \ram_block1a31~PORTBDATAOUT0 ;
wire \ram_block1a96~portadataout ;
wire \ram_block1a96~PORTBDATAOUT0 ;
wire \ram_block1a32~portadataout ;
wire \ram_block1a32~PORTBDATAOUT0 ;
wire \ram_block1a97~portadataout ;
wire \ram_block1a97~PORTBDATAOUT0 ;
wire \ram_block1a33~portadataout ;
wire \ram_block1a33~PORTBDATAOUT0 ;
wire \ram_block1a98~portadataout ;
wire \ram_block1a98~PORTBDATAOUT0 ;
wire \ram_block1a34~portadataout ;
wire \ram_block1a34~PORTBDATAOUT0 ;
wire \ram_block1a99~portadataout ;
wire \ram_block1a99~PORTBDATAOUT0 ;
wire \ram_block1a35~portadataout ;
wire \ram_block1a35~PORTBDATAOUT0 ;
wire \ram_block1a100~portadataout ;
wire \ram_block1a100~PORTBDATAOUT0 ;
wire \ram_block1a36~portadataout ;
wire \ram_block1a36~PORTBDATAOUT0 ;
wire \ram_block1a101~portadataout ;
wire \ram_block1a101~PORTBDATAOUT0 ;
wire \ram_block1a37~portadataout ;
wire \ram_block1a37~PORTBDATAOUT0 ;
wire \ram_block1a102~portadataout ;
wire \ram_block1a102~PORTBDATAOUT0 ;
wire \ram_block1a38~portadataout ;
wire \ram_block1a38~PORTBDATAOUT0 ;
wire \ram_block1a103~portadataout ;
wire \ram_block1a103~PORTBDATAOUT0 ;
wire \ram_block1a39~portadataout ;
wire \ram_block1a39~PORTBDATAOUT0 ;
wire \ram_block1a104~portadataout ;
wire \ram_block1a104~PORTBDATAOUT0 ;
wire \ram_block1a40~portadataout ;
wire \ram_block1a40~PORTBDATAOUT0 ;
wire \ram_block1a105~portadataout ;
wire \ram_block1a105~PORTBDATAOUT0 ;
wire \ram_block1a41~portadataout ;
wire \ram_block1a41~PORTBDATAOUT0 ;
wire \ram_block1a106~portadataout ;
wire \ram_block1a106~PORTBDATAOUT0 ;
wire \ram_block1a42~portadataout ;
wire \ram_block1a42~PORTBDATAOUT0 ;
wire \ram_block1a107~portadataout ;
wire \ram_block1a107~PORTBDATAOUT0 ;
wire \ram_block1a43~portadataout ;
wire \ram_block1a43~PORTBDATAOUT0 ;
wire \ram_block1a108~portadataout ;
wire \ram_block1a108~PORTBDATAOUT0 ;
wire \ram_block1a44~portadataout ;
wire \ram_block1a44~PORTBDATAOUT0 ;
wire \ram_block1a109~portadataout ;
wire \ram_block1a109~PORTBDATAOUT0 ;
wire \ram_block1a45~portadataout ;
wire \ram_block1a45~PORTBDATAOUT0 ;
wire \ram_block1a110~portadataout ;
wire \ram_block1a110~PORTBDATAOUT0 ;
wire \ram_block1a46~portadataout ;
wire \ram_block1a46~PORTBDATAOUT0 ;
wire \ram_block1a111~portadataout ;
wire \ram_block1a111~PORTBDATAOUT0 ;
wire \ram_block1a47~portadataout ;
wire \ram_block1a47~PORTBDATAOUT0 ;
wire \ram_block1a112~portadataout ;
wire \ram_block1a112~PORTBDATAOUT0 ;
wire \ram_block1a48~portadataout ;
wire \ram_block1a48~PORTBDATAOUT0 ;
wire \ram_block1a113~portadataout ;
wire \ram_block1a113~PORTBDATAOUT0 ;
wire \ram_block1a49~portadataout ;
wire \ram_block1a49~PORTBDATAOUT0 ;
wire \ram_block1a114~portadataout ;
wire \ram_block1a114~PORTBDATAOUT0 ;
wire \ram_block1a50~portadataout ;
wire \ram_block1a50~PORTBDATAOUT0 ;
wire \ram_block1a115~portadataout ;
wire \ram_block1a115~PORTBDATAOUT0 ;
wire \ram_block1a51~portadataout ;
wire \ram_block1a51~PORTBDATAOUT0 ;
wire \ram_block1a116~portadataout ;
wire \ram_block1a116~PORTBDATAOUT0 ;
wire \ram_block1a52~portadataout ;
wire \ram_block1a52~PORTBDATAOUT0 ;
wire \ram_block1a117~portadataout ;
wire \ram_block1a117~PORTBDATAOUT0 ;
wire \ram_block1a53~portadataout ;
wire \ram_block1a53~PORTBDATAOUT0 ;
wire \ram_block1a118~portadataout ;
wire \ram_block1a118~PORTBDATAOUT0 ;
wire \ram_block1a54~portadataout ;
wire \ram_block1a54~PORTBDATAOUT0 ;
wire \ram_block1a119~portadataout ;
wire \ram_block1a119~PORTBDATAOUT0 ;
wire \ram_block1a55~portadataout ;
wire \ram_block1a55~PORTBDATAOUT0 ;
wire \ram_block1a120~portadataout ;
wire \ram_block1a120~PORTBDATAOUT0 ;
wire \ram_block1a56~portadataout ;
wire \ram_block1a56~PORTBDATAOUT0 ;
wire \ram_block1a121~portadataout ;
wire \ram_block1a121~PORTBDATAOUT0 ;
wire \ram_block1a57~portadataout ;
wire \ram_block1a57~PORTBDATAOUT0 ;
wire \ram_block1a122~portadataout ;
wire \ram_block1a122~PORTBDATAOUT0 ;
wire \ram_block1a58~portadataout ;
wire \ram_block1a58~PORTBDATAOUT0 ;
wire \ram_block1a123~portadataout ;
wire \ram_block1a123~PORTBDATAOUT0 ;
wire \ram_block1a59~portadataout ;
wire \ram_block1a59~PORTBDATAOUT0 ;
wire \ram_block1a124~portadataout ;
wire \ram_block1a124~PORTBDATAOUT0 ;
wire \ram_block1a60~portadataout ;
wire \ram_block1a60~PORTBDATAOUT0 ;
wire \ram_block1a125~portadataout ;
wire \ram_block1a125~PORTBDATAOUT0 ;
wire \ram_block1a61~portadataout ;
wire \ram_block1a61~PORTBDATAOUT0 ;
wire \ram_block1a126~portadataout ;
wire \ram_block1a126~PORTBDATAOUT0 ;
wire \ram_block1a62~portadataout ;
wire \ram_block1a62~PORTBDATAOUT0 ;
wire \ram_block1a127~portadataout ;
wire \ram_block1a127~PORTBDATAOUT0 ;
wire \ram_block1a63~portadataout ;
wire \ram_block1a63~PORTBDATAOUT0 ;
wire \address_reg_a[0]~q ;
wire \address_reg_b[0]~q ;
wire \decode2|eq_node[1]~0_combout ;
wire \decode3|eq_node[1]~0_combout ;
wire \decode2|eq_node[0]~1_combout ;
wire \decode3|eq_node[0]~1_combout ;

wire [143:0] ram_block1a64_PORTADATAOUT_bus;
wire [143:0] ram_block1a64_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a65_PORTADATAOUT_bus;
wire [143:0] ram_block1a65_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a66_PORTADATAOUT_bus;
wire [143:0] ram_block1a66_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a67_PORTADATAOUT_bus;
wire [143:0] ram_block1a67_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a68_PORTADATAOUT_bus;
wire [143:0] ram_block1a68_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a69_PORTADATAOUT_bus;
wire [143:0] ram_block1a69_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a70_PORTADATAOUT_bus;
wire [143:0] ram_block1a70_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a71_PORTADATAOUT_bus;
wire [143:0] ram_block1a71_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a72_PORTADATAOUT_bus;
wire [143:0] ram_block1a72_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a73_PORTADATAOUT_bus;
wire [143:0] ram_block1a73_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a74_PORTADATAOUT_bus;
wire [143:0] ram_block1a74_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a75_PORTADATAOUT_bus;
wire [143:0] ram_block1a75_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a76_PORTADATAOUT_bus;
wire [143:0] ram_block1a76_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a77_PORTADATAOUT_bus;
wire [143:0] ram_block1a77_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a78_PORTADATAOUT_bus;
wire [143:0] ram_block1a78_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a79_PORTADATAOUT_bus;
wire [143:0] ram_block1a79_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a80_PORTADATAOUT_bus;
wire [143:0] ram_block1a80_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a81_PORTADATAOUT_bus;
wire [143:0] ram_block1a81_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a82_PORTADATAOUT_bus;
wire [143:0] ram_block1a82_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a83_PORTADATAOUT_bus;
wire [143:0] ram_block1a83_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a84_PORTADATAOUT_bus;
wire [143:0] ram_block1a84_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a85_PORTADATAOUT_bus;
wire [143:0] ram_block1a85_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a86_PORTADATAOUT_bus;
wire [143:0] ram_block1a86_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a87_PORTADATAOUT_bus;
wire [143:0] ram_block1a87_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a88_PORTADATAOUT_bus;
wire [143:0] ram_block1a88_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a89_PORTADATAOUT_bus;
wire [143:0] ram_block1a89_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a90_PORTADATAOUT_bus;
wire [143:0] ram_block1a90_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a91_PORTADATAOUT_bus;
wire [143:0] ram_block1a91_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a92_PORTADATAOUT_bus;
wire [143:0] ram_block1a92_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a93_PORTADATAOUT_bus;
wire [143:0] ram_block1a93_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a94_PORTADATAOUT_bus;
wire [143:0] ram_block1a94_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a95_PORTADATAOUT_bus;
wire [143:0] ram_block1a95_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a96_PORTADATAOUT_bus;
wire [143:0] ram_block1a96_PORTBDATAOUT_bus;
wire [143:0] ram_block1a32_PORTADATAOUT_bus;
wire [143:0] ram_block1a32_PORTBDATAOUT_bus;
wire [143:0] ram_block1a97_PORTADATAOUT_bus;
wire [143:0] ram_block1a97_PORTBDATAOUT_bus;
wire [143:0] ram_block1a33_PORTADATAOUT_bus;
wire [143:0] ram_block1a33_PORTBDATAOUT_bus;
wire [143:0] ram_block1a98_PORTADATAOUT_bus;
wire [143:0] ram_block1a98_PORTBDATAOUT_bus;
wire [143:0] ram_block1a34_PORTADATAOUT_bus;
wire [143:0] ram_block1a34_PORTBDATAOUT_bus;
wire [143:0] ram_block1a99_PORTADATAOUT_bus;
wire [143:0] ram_block1a99_PORTBDATAOUT_bus;
wire [143:0] ram_block1a35_PORTADATAOUT_bus;
wire [143:0] ram_block1a35_PORTBDATAOUT_bus;
wire [143:0] ram_block1a100_PORTADATAOUT_bus;
wire [143:0] ram_block1a100_PORTBDATAOUT_bus;
wire [143:0] ram_block1a36_PORTADATAOUT_bus;
wire [143:0] ram_block1a36_PORTBDATAOUT_bus;
wire [143:0] ram_block1a101_PORTADATAOUT_bus;
wire [143:0] ram_block1a101_PORTBDATAOUT_bus;
wire [143:0] ram_block1a37_PORTADATAOUT_bus;
wire [143:0] ram_block1a37_PORTBDATAOUT_bus;
wire [143:0] ram_block1a102_PORTADATAOUT_bus;
wire [143:0] ram_block1a102_PORTBDATAOUT_bus;
wire [143:0] ram_block1a38_PORTADATAOUT_bus;
wire [143:0] ram_block1a38_PORTBDATAOUT_bus;
wire [143:0] ram_block1a103_PORTADATAOUT_bus;
wire [143:0] ram_block1a103_PORTBDATAOUT_bus;
wire [143:0] ram_block1a39_PORTADATAOUT_bus;
wire [143:0] ram_block1a39_PORTBDATAOUT_bus;
wire [143:0] ram_block1a104_PORTADATAOUT_bus;
wire [143:0] ram_block1a104_PORTBDATAOUT_bus;
wire [143:0] ram_block1a40_PORTADATAOUT_bus;
wire [143:0] ram_block1a40_PORTBDATAOUT_bus;
wire [143:0] ram_block1a105_PORTADATAOUT_bus;
wire [143:0] ram_block1a105_PORTBDATAOUT_bus;
wire [143:0] ram_block1a41_PORTADATAOUT_bus;
wire [143:0] ram_block1a41_PORTBDATAOUT_bus;
wire [143:0] ram_block1a106_PORTADATAOUT_bus;
wire [143:0] ram_block1a106_PORTBDATAOUT_bus;
wire [143:0] ram_block1a42_PORTADATAOUT_bus;
wire [143:0] ram_block1a42_PORTBDATAOUT_bus;
wire [143:0] ram_block1a107_PORTADATAOUT_bus;
wire [143:0] ram_block1a107_PORTBDATAOUT_bus;
wire [143:0] ram_block1a43_PORTADATAOUT_bus;
wire [143:0] ram_block1a43_PORTBDATAOUT_bus;
wire [143:0] ram_block1a108_PORTADATAOUT_bus;
wire [143:0] ram_block1a108_PORTBDATAOUT_bus;
wire [143:0] ram_block1a44_PORTADATAOUT_bus;
wire [143:0] ram_block1a44_PORTBDATAOUT_bus;
wire [143:0] ram_block1a109_PORTADATAOUT_bus;
wire [143:0] ram_block1a109_PORTBDATAOUT_bus;
wire [143:0] ram_block1a45_PORTADATAOUT_bus;
wire [143:0] ram_block1a45_PORTBDATAOUT_bus;
wire [143:0] ram_block1a110_PORTADATAOUT_bus;
wire [143:0] ram_block1a110_PORTBDATAOUT_bus;
wire [143:0] ram_block1a46_PORTADATAOUT_bus;
wire [143:0] ram_block1a46_PORTBDATAOUT_bus;
wire [143:0] ram_block1a111_PORTADATAOUT_bus;
wire [143:0] ram_block1a111_PORTBDATAOUT_bus;
wire [143:0] ram_block1a47_PORTADATAOUT_bus;
wire [143:0] ram_block1a47_PORTBDATAOUT_bus;
wire [143:0] ram_block1a112_PORTADATAOUT_bus;
wire [143:0] ram_block1a112_PORTBDATAOUT_bus;
wire [143:0] ram_block1a48_PORTADATAOUT_bus;
wire [143:0] ram_block1a48_PORTBDATAOUT_bus;
wire [143:0] ram_block1a113_PORTADATAOUT_bus;
wire [143:0] ram_block1a113_PORTBDATAOUT_bus;
wire [143:0] ram_block1a49_PORTADATAOUT_bus;
wire [143:0] ram_block1a49_PORTBDATAOUT_bus;
wire [143:0] ram_block1a114_PORTADATAOUT_bus;
wire [143:0] ram_block1a114_PORTBDATAOUT_bus;
wire [143:0] ram_block1a50_PORTADATAOUT_bus;
wire [143:0] ram_block1a50_PORTBDATAOUT_bus;
wire [143:0] ram_block1a115_PORTADATAOUT_bus;
wire [143:0] ram_block1a115_PORTBDATAOUT_bus;
wire [143:0] ram_block1a51_PORTADATAOUT_bus;
wire [143:0] ram_block1a51_PORTBDATAOUT_bus;
wire [143:0] ram_block1a116_PORTADATAOUT_bus;
wire [143:0] ram_block1a116_PORTBDATAOUT_bus;
wire [143:0] ram_block1a52_PORTADATAOUT_bus;
wire [143:0] ram_block1a52_PORTBDATAOUT_bus;
wire [143:0] ram_block1a117_PORTADATAOUT_bus;
wire [143:0] ram_block1a117_PORTBDATAOUT_bus;
wire [143:0] ram_block1a53_PORTADATAOUT_bus;
wire [143:0] ram_block1a53_PORTBDATAOUT_bus;
wire [143:0] ram_block1a118_PORTADATAOUT_bus;
wire [143:0] ram_block1a118_PORTBDATAOUT_bus;
wire [143:0] ram_block1a54_PORTADATAOUT_bus;
wire [143:0] ram_block1a54_PORTBDATAOUT_bus;
wire [143:0] ram_block1a119_PORTADATAOUT_bus;
wire [143:0] ram_block1a119_PORTBDATAOUT_bus;
wire [143:0] ram_block1a55_PORTADATAOUT_bus;
wire [143:0] ram_block1a55_PORTBDATAOUT_bus;
wire [143:0] ram_block1a120_PORTADATAOUT_bus;
wire [143:0] ram_block1a120_PORTBDATAOUT_bus;
wire [143:0] ram_block1a56_PORTADATAOUT_bus;
wire [143:0] ram_block1a56_PORTBDATAOUT_bus;
wire [143:0] ram_block1a121_PORTADATAOUT_bus;
wire [143:0] ram_block1a121_PORTBDATAOUT_bus;
wire [143:0] ram_block1a57_PORTADATAOUT_bus;
wire [143:0] ram_block1a57_PORTBDATAOUT_bus;
wire [143:0] ram_block1a122_PORTADATAOUT_bus;
wire [143:0] ram_block1a122_PORTBDATAOUT_bus;
wire [143:0] ram_block1a58_PORTADATAOUT_bus;
wire [143:0] ram_block1a58_PORTBDATAOUT_bus;
wire [143:0] ram_block1a123_PORTADATAOUT_bus;
wire [143:0] ram_block1a123_PORTBDATAOUT_bus;
wire [143:0] ram_block1a59_PORTADATAOUT_bus;
wire [143:0] ram_block1a59_PORTBDATAOUT_bus;
wire [143:0] ram_block1a124_PORTADATAOUT_bus;
wire [143:0] ram_block1a124_PORTBDATAOUT_bus;
wire [143:0] ram_block1a60_PORTADATAOUT_bus;
wire [143:0] ram_block1a60_PORTBDATAOUT_bus;
wire [143:0] ram_block1a125_PORTADATAOUT_bus;
wire [143:0] ram_block1a125_PORTBDATAOUT_bus;
wire [143:0] ram_block1a61_PORTADATAOUT_bus;
wire [143:0] ram_block1a61_PORTBDATAOUT_bus;
wire [143:0] ram_block1a126_PORTADATAOUT_bus;
wire [143:0] ram_block1a126_PORTBDATAOUT_bus;
wire [143:0] ram_block1a62_PORTADATAOUT_bus;
wire [143:0] ram_block1a62_PORTBDATAOUT_bus;
wire [143:0] ram_block1a127_PORTADATAOUT_bus;
wire [143:0] ram_block1a127_PORTBDATAOUT_bus;
wire [143:0] ram_block1a63_PORTADATAOUT_bus;
wire [143:0] ram_block1a63_PORTBDATAOUT_bus;

assign \ram_block1a64~portadataout  = ram_block1a64_PORTADATAOUT_bus[0];

assign \ram_block1a64~PORTBDATAOUT0  = ram_block1a64_PORTBDATAOUT_bus[0];

assign \ram_block1a0~portadataout  = ram_block1a0_PORTADATAOUT_bus[0];

assign \ram_block1a0~PORTBDATAOUT0  = ram_block1a0_PORTBDATAOUT_bus[0];

assign \ram_block1a65~portadataout  = ram_block1a65_PORTADATAOUT_bus[0];

assign \ram_block1a65~PORTBDATAOUT0  = ram_block1a65_PORTBDATAOUT_bus[0];

assign \ram_block1a1~portadataout  = ram_block1a1_PORTADATAOUT_bus[0];

assign \ram_block1a1~PORTBDATAOUT0  = ram_block1a1_PORTBDATAOUT_bus[0];

assign \ram_block1a66~portadataout  = ram_block1a66_PORTADATAOUT_bus[0];

assign \ram_block1a66~PORTBDATAOUT0  = ram_block1a66_PORTBDATAOUT_bus[0];

assign \ram_block1a2~portadataout  = ram_block1a2_PORTADATAOUT_bus[0];

assign \ram_block1a2~PORTBDATAOUT0  = ram_block1a2_PORTBDATAOUT_bus[0];

assign \ram_block1a67~portadataout  = ram_block1a67_PORTADATAOUT_bus[0];

assign \ram_block1a67~PORTBDATAOUT0  = ram_block1a67_PORTBDATAOUT_bus[0];

assign \ram_block1a3~portadataout  = ram_block1a3_PORTADATAOUT_bus[0];

assign \ram_block1a3~PORTBDATAOUT0  = ram_block1a3_PORTBDATAOUT_bus[0];

assign \ram_block1a68~portadataout  = ram_block1a68_PORTADATAOUT_bus[0];

assign \ram_block1a68~PORTBDATAOUT0  = ram_block1a68_PORTBDATAOUT_bus[0];

assign \ram_block1a4~portadataout  = ram_block1a4_PORTADATAOUT_bus[0];

assign \ram_block1a4~PORTBDATAOUT0  = ram_block1a4_PORTBDATAOUT_bus[0];

assign \ram_block1a69~portadataout  = ram_block1a69_PORTADATAOUT_bus[0];

assign \ram_block1a69~PORTBDATAOUT0  = ram_block1a69_PORTBDATAOUT_bus[0];

assign \ram_block1a5~portadataout  = ram_block1a5_PORTADATAOUT_bus[0];

assign \ram_block1a5~PORTBDATAOUT0  = ram_block1a5_PORTBDATAOUT_bus[0];

assign \ram_block1a70~portadataout  = ram_block1a70_PORTADATAOUT_bus[0];

assign \ram_block1a70~PORTBDATAOUT0  = ram_block1a70_PORTBDATAOUT_bus[0];

assign \ram_block1a6~portadataout  = ram_block1a6_PORTADATAOUT_bus[0];

assign \ram_block1a6~PORTBDATAOUT0  = ram_block1a6_PORTBDATAOUT_bus[0];

assign \ram_block1a71~portadataout  = ram_block1a71_PORTADATAOUT_bus[0];

assign \ram_block1a71~PORTBDATAOUT0  = ram_block1a71_PORTBDATAOUT_bus[0];

assign \ram_block1a7~portadataout  = ram_block1a7_PORTADATAOUT_bus[0];

assign \ram_block1a7~PORTBDATAOUT0  = ram_block1a7_PORTBDATAOUT_bus[0];

assign \ram_block1a72~portadataout  = ram_block1a72_PORTADATAOUT_bus[0];

assign \ram_block1a72~PORTBDATAOUT0  = ram_block1a72_PORTBDATAOUT_bus[0];

assign \ram_block1a8~portadataout  = ram_block1a8_PORTADATAOUT_bus[0];

assign \ram_block1a8~PORTBDATAOUT0  = ram_block1a8_PORTBDATAOUT_bus[0];

assign \ram_block1a73~portadataout  = ram_block1a73_PORTADATAOUT_bus[0];

assign \ram_block1a73~PORTBDATAOUT0  = ram_block1a73_PORTBDATAOUT_bus[0];

assign \ram_block1a9~portadataout  = ram_block1a9_PORTADATAOUT_bus[0];

assign \ram_block1a9~PORTBDATAOUT0  = ram_block1a9_PORTBDATAOUT_bus[0];

assign \ram_block1a74~portadataout  = ram_block1a74_PORTADATAOUT_bus[0];

assign \ram_block1a74~PORTBDATAOUT0  = ram_block1a74_PORTBDATAOUT_bus[0];

assign \ram_block1a10~portadataout  = ram_block1a10_PORTADATAOUT_bus[0];

assign \ram_block1a10~PORTBDATAOUT0  = ram_block1a10_PORTBDATAOUT_bus[0];

assign \ram_block1a75~portadataout  = ram_block1a75_PORTADATAOUT_bus[0];

assign \ram_block1a75~PORTBDATAOUT0  = ram_block1a75_PORTBDATAOUT_bus[0];

assign \ram_block1a11~portadataout  = ram_block1a11_PORTADATAOUT_bus[0];

assign \ram_block1a11~PORTBDATAOUT0  = ram_block1a11_PORTBDATAOUT_bus[0];

assign \ram_block1a76~portadataout  = ram_block1a76_PORTADATAOUT_bus[0];

assign \ram_block1a76~PORTBDATAOUT0  = ram_block1a76_PORTBDATAOUT_bus[0];

assign \ram_block1a12~portadataout  = ram_block1a12_PORTADATAOUT_bus[0];

assign \ram_block1a12~PORTBDATAOUT0  = ram_block1a12_PORTBDATAOUT_bus[0];

assign \ram_block1a77~portadataout  = ram_block1a77_PORTADATAOUT_bus[0];

assign \ram_block1a77~PORTBDATAOUT0  = ram_block1a77_PORTBDATAOUT_bus[0];

assign \ram_block1a13~portadataout  = ram_block1a13_PORTADATAOUT_bus[0];

assign \ram_block1a13~PORTBDATAOUT0  = ram_block1a13_PORTBDATAOUT_bus[0];

assign \ram_block1a78~portadataout  = ram_block1a78_PORTADATAOUT_bus[0];

assign \ram_block1a78~PORTBDATAOUT0  = ram_block1a78_PORTBDATAOUT_bus[0];

assign \ram_block1a14~portadataout  = ram_block1a14_PORTADATAOUT_bus[0];

assign \ram_block1a14~PORTBDATAOUT0  = ram_block1a14_PORTBDATAOUT_bus[0];

assign \ram_block1a79~portadataout  = ram_block1a79_PORTADATAOUT_bus[0];

assign \ram_block1a79~PORTBDATAOUT0  = ram_block1a79_PORTBDATAOUT_bus[0];

assign \ram_block1a15~portadataout  = ram_block1a15_PORTADATAOUT_bus[0];

assign \ram_block1a15~PORTBDATAOUT0  = ram_block1a15_PORTBDATAOUT_bus[0];

assign \ram_block1a80~portadataout  = ram_block1a80_PORTADATAOUT_bus[0];

assign \ram_block1a80~PORTBDATAOUT0  = ram_block1a80_PORTBDATAOUT_bus[0];

assign \ram_block1a16~portadataout  = ram_block1a16_PORTADATAOUT_bus[0];

assign \ram_block1a16~PORTBDATAOUT0  = ram_block1a16_PORTBDATAOUT_bus[0];

assign \ram_block1a81~portadataout  = ram_block1a81_PORTADATAOUT_bus[0];

assign \ram_block1a81~PORTBDATAOUT0  = ram_block1a81_PORTBDATAOUT_bus[0];

assign \ram_block1a17~portadataout  = ram_block1a17_PORTADATAOUT_bus[0];

assign \ram_block1a17~PORTBDATAOUT0  = ram_block1a17_PORTBDATAOUT_bus[0];

assign \ram_block1a82~portadataout  = ram_block1a82_PORTADATAOUT_bus[0];

assign \ram_block1a82~PORTBDATAOUT0  = ram_block1a82_PORTBDATAOUT_bus[0];

assign \ram_block1a18~portadataout  = ram_block1a18_PORTADATAOUT_bus[0];

assign \ram_block1a18~PORTBDATAOUT0  = ram_block1a18_PORTBDATAOUT_bus[0];

assign \ram_block1a83~portadataout  = ram_block1a83_PORTADATAOUT_bus[0];

assign \ram_block1a83~PORTBDATAOUT0  = ram_block1a83_PORTBDATAOUT_bus[0];

assign \ram_block1a19~portadataout  = ram_block1a19_PORTADATAOUT_bus[0];

assign \ram_block1a19~PORTBDATAOUT0  = ram_block1a19_PORTBDATAOUT_bus[0];

assign \ram_block1a84~portadataout  = ram_block1a84_PORTADATAOUT_bus[0];

assign \ram_block1a84~PORTBDATAOUT0  = ram_block1a84_PORTBDATAOUT_bus[0];

assign \ram_block1a20~portadataout  = ram_block1a20_PORTADATAOUT_bus[0];

assign \ram_block1a20~PORTBDATAOUT0  = ram_block1a20_PORTBDATAOUT_bus[0];

assign \ram_block1a85~portadataout  = ram_block1a85_PORTADATAOUT_bus[0];

assign \ram_block1a85~PORTBDATAOUT0  = ram_block1a85_PORTBDATAOUT_bus[0];

assign \ram_block1a21~portadataout  = ram_block1a21_PORTADATAOUT_bus[0];

assign \ram_block1a21~PORTBDATAOUT0  = ram_block1a21_PORTBDATAOUT_bus[0];

assign \ram_block1a86~portadataout  = ram_block1a86_PORTADATAOUT_bus[0];

assign \ram_block1a86~PORTBDATAOUT0  = ram_block1a86_PORTBDATAOUT_bus[0];

assign \ram_block1a22~portadataout  = ram_block1a22_PORTADATAOUT_bus[0];

assign \ram_block1a22~PORTBDATAOUT0  = ram_block1a22_PORTBDATAOUT_bus[0];

assign \ram_block1a87~portadataout  = ram_block1a87_PORTADATAOUT_bus[0];

assign \ram_block1a87~PORTBDATAOUT0  = ram_block1a87_PORTBDATAOUT_bus[0];

assign \ram_block1a23~portadataout  = ram_block1a23_PORTADATAOUT_bus[0];

assign \ram_block1a23~PORTBDATAOUT0  = ram_block1a23_PORTBDATAOUT_bus[0];

assign \ram_block1a88~portadataout  = ram_block1a88_PORTADATAOUT_bus[0];

assign \ram_block1a88~PORTBDATAOUT0  = ram_block1a88_PORTBDATAOUT_bus[0];

assign \ram_block1a24~portadataout  = ram_block1a24_PORTADATAOUT_bus[0];

assign \ram_block1a24~PORTBDATAOUT0  = ram_block1a24_PORTBDATAOUT_bus[0];

assign \ram_block1a89~portadataout  = ram_block1a89_PORTADATAOUT_bus[0];

assign \ram_block1a89~PORTBDATAOUT0  = ram_block1a89_PORTBDATAOUT_bus[0];

assign \ram_block1a25~portadataout  = ram_block1a25_PORTADATAOUT_bus[0];

assign \ram_block1a25~PORTBDATAOUT0  = ram_block1a25_PORTBDATAOUT_bus[0];

assign \ram_block1a90~portadataout  = ram_block1a90_PORTADATAOUT_bus[0];

assign \ram_block1a90~PORTBDATAOUT0  = ram_block1a90_PORTBDATAOUT_bus[0];

assign \ram_block1a26~portadataout  = ram_block1a26_PORTADATAOUT_bus[0];

assign \ram_block1a26~PORTBDATAOUT0  = ram_block1a26_PORTBDATAOUT_bus[0];

assign \ram_block1a91~portadataout  = ram_block1a91_PORTADATAOUT_bus[0];

assign \ram_block1a91~PORTBDATAOUT0  = ram_block1a91_PORTBDATAOUT_bus[0];

assign \ram_block1a27~portadataout  = ram_block1a27_PORTADATAOUT_bus[0];

assign \ram_block1a27~PORTBDATAOUT0  = ram_block1a27_PORTBDATAOUT_bus[0];

assign \ram_block1a92~portadataout  = ram_block1a92_PORTADATAOUT_bus[0];

assign \ram_block1a92~PORTBDATAOUT0  = ram_block1a92_PORTBDATAOUT_bus[0];

assign \ram_block1a28~portadataout  = ram_block1a28_PORTADATAOUT_bus[0];

assign \ram_block1a28~PORTBDATAOUT0  = ram_block1a28_PORTBDATAOUT_bus[0];

assign \ram_block1a93~portadataout  = ram_block1a93_PORTADATAOUT_bus[0];

assign \ram_block1a93~PORTBDATAOUT0  = ram_block1a93_PORTBDATAOUT_bus[0];

assign \ram_block1a29~portadataout  = ram_block1a29_PORTADATAOUT_bus[0];

assign \ram_block1a29~PORTBDATAOUT0  = ram_block1a29_PORTBDATAOUT_bus[0];

assign \ram_block1a94~portadataout  = ram_block1a94_PORTADATAOUT_bus[0];

assign \ram_block1a94~PORTBDATAOUT0  = ram_block1a94_PORTBDATAOUT_bus[0];

assign \ram_block1a30~portadataout  = ram_block1a30_PORTADATAOUT_bus[0];

assign \ram_block1a30~PORTBDATAOUT0  = ram_block1a30_PORTBDATAOUT_bus[0];

assign \ram_block1a95~portadataout  = ram_block1a95_PORTADATAOUT_bus[0];

assign \ram_block1a95~PORTBDATAOUT0  = ram_block1a95_PORTBDATAOUT_bus[0];

assign \ram_block1a31~portadataout  = ram_block1a31_PORTADATAOUT_bus[0];

assign \ram_block1a31~PORTBDATAOUT0  = ram_block1a31_PORTBDATAOUT_bus[0];

assign \ram_block1a96~portadataout  = ram_block1a96_PORTADATAOUT_bus[0];

assign \ram_block1a96~PORTBDATAOUT0  = ram_block1a96_PORTBDATAOUT_bus[0];

assign \ram_block1a32~portadataout  = ram_block1a32_PORTADATAOUT_bus[0];

assign \ram_block1a32~PORTBDATAOUT0  = ram_block1a32_PORTBDATAOUT_bus[0];

assign \ram_block1a97~portadataout  = ram_block1a97_PORTADATAOUT_bus[0];

assign \ram_block1a97~PORTBDATAOUT0  = ram_block1a97_PORTBDATAOUT_bus[0];

assign \ram_block1a33~portadataout  = ram_block1a33_PORTADATAOUT_bus[0];

assign \ram_block1a33~PORTBDATAOUT0  = ram_block1a33_PORTBDATAOUT_bus[0];

assign \ram_block1a98~portadataout  = ram_block1a98_PORTADATAOUT_bus[0];

assign \ram_block1a98~PORTBDATAOUT0  = ram_block1a98_PORTBDATAOUT_bus[0];

assign \ram_block1a34~portadataout  = ram_block1a34_PORTADATAOUT_bus[0];

assign \ram_block1a34~PORTBDATAOUT0  = ram_block1a34_PORTBDATAOUT_bus[0];

assign \ram_block1a99~portadataout  = ram_block1a99_PORTADATAOUT_bus[0];

assign \ram_block1a99~PORTBDATAOUT0  = ram_block1a99_PORTBDATAOUT_bus[0];

assign \ram_block1a35~portadataout  = ram_block1a35_PORTADATAOUT_bus[0];

assign \ram_block1a35~PORTBDATAOUT0  = ram_block1a35_PORTBDATAOUT_bus[0];

assign \ram_block1a100~portadataout  = ram_block1a100_PORTADATAOUT_bus[0];

assign \ram_block1a100~PORTBDATAOUT0  = ram_block1a100_PORTBDATAOUT_bus[0];

assign \ram_block1a36~portadataout  = ram_block1a36_PORTADATAOUT_bus[0];

assign \ram_block1a36~PORTBDATAOUT0  = ram_block1a36_PORTBDATAOUT_bus[0];

assign \ram_block1a101~portadataout  = ram_block1a101_PORTADATAOUT_bus[0];

assign \ram_block1a101~PORTBDATAOUT0  = ram_block1a101_PORTBDATAOUT_bus[0];

assign \ram_block1a37~portadataout  = ram_block1a37_PORTADATAOUT_bus[0];

assign \ram_block1a37~PORTBDATAOUT0  = ram_block1a37_PORTBDATAOUT_bus[0];

assign \ram_block1a102~portadataout  = ram_block1a102_PORTADATAOUT_bus[0];

assign \ram_block1a102~PORTBDATAOUT0  = ram_block1a102_PORTBDATAOUT_bus[0];

assign \ram_block1a38~portadataout  = ram_block1a38_PORTADATAOUT_bus[0];

assign \ram_block1a38~PORTBDATAOUT0  = ram_block1a38_PORTBDATAOUT_bus[0];

assign \ram_block1a103~portadataout  = ram_block1a103_PORTADATAOUT_bus[0];

assign \ram_block1a103~PORTBDATAOUT0  = ram_block1a103_PORTBDATAOUT_bus[0];

assign \ram_block1a39~portadataout  = ram_block1a39_PORTADATAOUT_bus[0];

assign \ram_block1a39~PORTBDATAOUT0  = ram_block1a39_PORTBDATAOUT_bus[0];

assign \ram_block1a104~portadataout  = ram_block1a104_PORTADATAOUT_bus[0];

assign \ram_block1a104~PORTBDATAOUT0  = ram_block1a104_PORTBDATAOUT_bus[0];

assign \ram_block1a40~portadataout  = ram_block1a40_PORTADATAOUT_bus[0];

assign \ram_block1a40~PORTBDATAOUT0  = ram_block1a40_PORTBDATAOUT_bus[0];

assign \ram_block1a105~portadataout  = ram_block1a105_PORTADATAOUT_bus[0];

assign \ram_block1a105~PORTBDATAOUT0  = ram_block1a105_PORTBDATAOUT_bus[0];

assign \ram_block1a41~portadataout  = ram_block1a41_PORTADATAOUT_bus[0];

assign \ram_block1a41~PORTBDATAOUT0  = ram_block1a41_PORTBDATAOUT_bus[0];

assign \ram_block1a106~portadataout  = ram_block1a106_PORTADATAOUT_bus[0];

assign \ram_block1a106~PORTBDATAOUT0  = ram_block1a106_PORTBDATAOUT_bus[0];

assign \ram_block1a42~portadataout  = ram_block1a42_PORTADATAOUT_bus[0];

assign \ram_block1a42~PORTBDATAOUT0  = ram_block1a42_PORTBDATAOUT_bus[0];

assign \ram_block1a107~portadataout  = ram_block1a107_PORTADATAOUT_bus[0];

assign \ram_block1a107~PORTBDATAOUT0  = ram_block1a107_PORTBDATAOUT_bus[0];

assign \ram_block1a43~portadataout  = ram_block1a43_PORTADATAOUT_bus[0];

assign \ram_block1a43~PORTBDATAOUT0  = ram_block1a43_PORTBDATAOUT_bus[0];

assign \ram_block1a108~portadataout  = ram_block1a108_PORTADATAOUT_bus[0];

assign \ram_block1a108~PORTBDATAOUT0  = ram_block1a108_PORTBDATAOUT_bus[0];

assign \ram_block1a44~portadataout  = ram_block1a44_PORTADATAOUT_bus[0];

assign \ram_block1a44~PORTBDATAOUT0  = ram_block1a44_PORTBDATAOUT_bus[0];

assign \ram_block1a109~portadataout  = ram_block1a109_PORTADATAOUT_bus[0];

assign \ram_block1a109~PORTBDATAOUT0  = ram_block1a109_PORTBDATAOUT_bus[0];

assign \ram_block1a45~portadataout  = ram_block1a45_PORTADATAOUT_bus[0];

assign \ram_block1a45~PORTBDATAOUT0  = ram_block1a45_PORTBDATAOUT_bus[0];

assign \ram_block1a110~portadataout  = ram_block1a110_PORTADATAOUT_bus[0];

assign \ram_block1a110~PORTBDATAOUT0  = ram_block1a110_PORTBDATAOUT_bus[0];

assign \ram_block1a46~portadataout  = ram_block1a46_PORTADATAOUT_bus[0];

assign \ram_block1a46~PORTBDATAOUT0  = ram_block1a46_PORTBDATAOUT_bus[0];

assign \ram_block1a111~portadataout  = ram_block1a111_PORTADATAOUT_bus[0];

assign \ram_block1a111~PORTBDATAOUT0  = ram_block1a111_PORTBDATAOUT_bus[0];

assign \ram_block1a47~portadataout  = ram_block1a47_PORTADATAOUT_bus[0];

assign \ram_block1a47~PORTBDATAOUT0  = ram_block1a47_PORTBDATAOUT_bus[0];

assign \ram_block1a112~portadataout  = ram_block1a112_PORTADATAOUT_bus[0];

assign \ram_block1a112~PORTBDATAOUT0  = ram_block1a112_PORTBDATAOUT_bus[0];

assign \ram_block1a48~portadataout  = ram_block1a48_PORTADATAOUT_bus[0];

assign \ram_block1a48~PORTBDATAOUT0  = ram_block1a48_PORTBDATAOUT_bus[0];

assign \ram_block1a113~portadataout  = ram_block1a113_PORTADATAOUT_bus[0];

assign \ram_block1a113~PORTBDATAOUT0  = ram_block1a113_PORTBDATAOUT_bus[0];

assign \ram_block1a49~portadataout  = ram_block1a49_PORTADATAOUT_bus[0];

assign \ram_block1a49~PORTBDATAOUT0  = ram_block1a49_PORTBDATAOUT_bus[0];

assign \ram_block1a114~portadataout  = ram_block1a114_PORTADATAOUT_bus[0];

assign \ram_block1a114~PORTBDATAOUT0  = ram_block1a114_PORTBDATAOUT_bus[0];

assign \ram_block1a50~portadataout  = ram_block1a50_PORTADATAOUT_bus[0];

assign \ram_block1a50~PORTBDATAOUT0  = ram_block1a50_PORTBDATAOUT_bus[0];

assign \ram_block1a115~portadataout  = ram_block1a115_PORTADATAOUT_bus[0];

assign \ram_block1a115~PORTBDATAOUT0  = ram_block1a115_PORTBDATAOUT_bus[0];

assign \ram_block1a51~portadataout  = ram_block1a51_PORTADATAOUT_bus[0];

assign \ram_block1a51~PORTBDATAOUT0  = ram_block1a51_PORTBDATAOUT_bus[0];

assign \ram_block1a116~portadataout  = ram_block1a116_PORTADATAOUT_bus[0];

assign \ram_block1a116~PORTBDATAOUT0  = ram_block1a116_PORTBDATAOUT_bus[0];

assign \ram_block1a52~portadataout  = ram_block1a52_PORTADATAOUT_bus[0];

assign \ram_block1a52~PORTBDATAOUT0  = ram_block1a52_PORTBDATAOUT_bus[0];

assign \ram_block1a117~portadataout  = ram_block1a117_PORTADATAOUT_bus[0];

assign \ram_block1a117~PORTBDATAOUT0  = ram_block1a117_PORTBDATAOUT_bus[0];

assign \ram_block1a53~portadataout  = ram_block1a53_PORTADATAOUT_bus[0];

assign \ram_block1a53~PORTBDATAOUT0  = ram_block1a53_PORTBDATAOUT_bus[0];

assign \ram_block1a118~portadataout  = ram_block1a118_PORTADATAOUT_bus[0];

assign \ram_block1a118~PORTBDATAOUT0  = ram_block1a118_PORTBDATAOUT_bus[0];

assign \ram_block1a54~portadataout  = ram_block1a54_PORTADATAOUT_bus[0];

assign \ram_block1a54~PORTBDATAOUT0  = ram_block1a54_PORTBDATAOUT_bus[0];

assign \ram_block1a119~portadataout  = ram_block1a119_PORTADATAOUT_bus[0];

assign \ram_block1a119~PORTBDATAOUT0  = ram_block1a119_PORTBDATAOUT_bus[0];

assign \ram_block1a55~portadataout  = ram_block1a55_PORTADATAOUT_bus[0];

assign \ram_block1a55~PORTBDATAOUT0  = ram_block1a55_PORTBDATAOUT_bus[0];

assign \ram_block1a120~portadataout  = ram_block1a120_PORTADATAOUT_bus[0];

assign \ram_block1a120~PORTBDATAOUT0  = ram_block1a120_PORTBDATAOUT_bus[0];

assign \ram_block1a56~portadataout  = ram_block1a56_PORTADATAOUT_bus[0];

assign \ram_block1a56~PORTBDATAOUT0  = ram_block1a56_PORTBDATAOUT_bus[0];

assign \ram_block1a121~portadataout  = ram_block1a121_PORTADATAOUT_bus[0];

assign \ram_block1a121~PORTBDATAOUT0  = ram_block1a121_PORTBDATAOUT_bus[0];

assign \ram_block1a57~portadataout  = ram_block1a57_PORTADATAOUT_bus[0];

assign \ram_block1a57~PORTBDATAOUT0  = ram_block1a57_PORTBDATAOUT_bus[0];

assign \ram_block1a122~portadataout  = ram_block1a122_PORTADATAOUT_bus[0];

assign \ram_block1a122~PORTBDATAOUT0  = ram_block1a122_PORTBDATAOUT_bus[0];

assign \ram_block1a58~portadataout  = ram_block1a58_PORTADATAOUT_bus[0];

assign \ram_block1a58~PORTBDATAOUT0  = ram_block1a58_PORTBDATAOUT_bus[0];

assign \ram_block1a123~portadataout  = ram_block1a123_PORTADATAOUT_bus[0];

assign \ram_block1a123~PORTBDATAOUT0  = ram_block1a123_PORTBDATAOUT_bus[0];

assign \ram_block1a59~portadataout  = ram_block1a59_PORTADATAOUT_bus[0];

assign \ram_block1a59~PORTBDATAOUT0  = ram_block1a59_PORTBDATAOUT_bus[0];

assign \ram_block1a124~portadataout  = ram_block1a124_PORTADATAOUT_bus[0];

assign \ram_block1a124~PORTBDATAOUT0  = ram_block1a124_PORTBDATAOUT_bus[0];

assign \ram_block1a60~portadataout  = ram_block1a60_PORTADATAOUT_bus[0];

assign \ram_block1a60~PORTBDATAOUT0  = ram_block1a60_PORTBDATAOUT_bus[0];

assign \ram_block1a125~portadataout  = ram_block1a125_PORTADATAOUT_bus[0];

assign \ram_block1a125~PORTBDATAOUT0  = ram_block1a125_PORTBDATAOUT_bus[0];

assign \ram_block1a61~portadataout  = ram_block1a61_PORTADATAOUT_bus[0];

assign \ram_block1a61~PORTBDATAOUT0  = ram_block1a61_PORTBDATAOUT_bus[0];

assign \ram_block1a126~portadataout  = ram_block1a126_PORTADATAOUT_bus[0];

assign \ram_block1a126~PORTBDATAOUT0  = ram_block1a126_PORTBDATAOUT_bus[0];

assign \ram_block1a62~portadataout  = ram_block1a62_PORTADATAOUT_bus[0];

assign \ram_block1a62~PORTBDATAOUT0  = ram_block1a62_PORTBDATAOUT_bus[0];

assign \ram_block1a127~portadataout  = ram_block1a127_PORTADATAOUT_bus[0];

assign \ram_block1a127~PORTBDATAOUT0  = ram_block1a127_PORTBDATAOUT_bus[0];

assign \ram_block1a63~portadataout  = ram_block1a63_PORTADATAOUT_bus[0];

assign \ram_block1a63~PORTBDATAOUT0  = ram_block1a63_PORTBDATAOUT_bus[0];

qtestpd_mux_fsb_1 mux5(
	.ram_block1a64(\ram_block1a64~PORTBDATAOUT0 ),
	.ram_block1a0(\ram_block1a0~PORTBDATAOUT0 ),
	.ram_block1a65(\ram_block1a65~PORTBDATAOUT0 ),
	.ram_block1a1(\ram_block1a1~PORTBDATAOUT0 ),
	.ram_block1a66(\ram_block1a66~PORTBDATAOUT0 ),
	.ram_block1a2(\ram_block1a2~PORTBDATAOUT0 ),
	.ram_block1a67(\ram_block1a67~PORTBDATAOUT0 ),
	.ram_block1a3(\ram_block1a3~PORTBDATAOUT0 ),
	.ram_block1a68(\ram_block1a68~PORTBDATAOUT0 ),
	.ram_block1a4(\ram_block1a4~PORTBDATAOUT0 ),
	.ram_block1a69(\ram_block1a69~PORTBDATAOUT0 ),
	.ram_block1a5(\ram_block1a5~PORTBDATAOUT0 ),
	.ram_block1a70(\ram_block1a70~PORTBDATAOUT0 ),
	.ram_block1a6(\ram_block1a6~PORTBDATAOUT0 ),
	.ram_block1a71(\ram_block1a71~PORTBDATAOUT0 ),
	.ram_block1a7(\ram_block1a7~PORTBDATAOUT0 ),
	.ram_block1a72(\ram_block1a72~PORTBDATAOUT0 ),
	.ram_block1a8(\ram_block1a8~PORTBDATAOUT0 ),
	.ram_block1a73(\ram_block1a73~PORTBDATAOUT0 ),
	.ram_block1a9(\ram_block1a9~PORTBDATAOUT0 ),
	.ram_block1a74(\ram_block1a74~PORTBDATAOUT0 ),
	.ram_block1a10(\ram_block1a10~PORTBDATAOUT0 ),
	.ram_block1a75(\ram_block1a75~PORTBDATAOUT0 ),
	.ram_block1a11(\ram_block1a11~PORTBDATAOUT0 ),
	.ram_block1a76(\ram_block1a76~PORTBDATAOUT0 ),
	.ram_block1a12(\ram_block1a12~PORTBDATAOUT0 ),
	.ram_block1a77(\ram_block1a77~PORTBDATAOUT0 ),
	.ram_block1a13(\ram_block1a13~PORTBDATAOUT0 ),
	.ram_block1a78(\ram_block1a78~PORTBDATAOUT0 ),
	.ram_block1a14(\ram_block1a14~PORTBDATAOUT0 ),
	.ram_block1a79(\ram_block1a79~PORTBDATAOUT0 ),
	.ram_block1a15(\ram_block1a15~PORTBDATAOUT0 ),
	.ram_block1a80(\ram_block1a80~PORTBDATAOUT0 ),
	.ram_block1a16(\ram_block1a16~PORTBDATAOUT0 ),
	.ram_block1a81(\ram_block1a81~PORTBDATAOUT0 ),
	.ram_block1a17(\ram_block1a17~PORTBDATAOUT0 ),
	.ram_block1a82(\ram_block1a82~PORTBDATAOUT0 ),
	.ram_block1a18(\ram_block1a18~PORTBDATAOUT0 ),
	.ram_block1a83(\ram_block1a83~PORTBDATAOUT0 ),
	.ram_block1a19(\ram_block1a19~PORTBDATAOUT0 ),
	.ram_block1a84(\ram_block1a84~PORTBDATAOUT0 ),
	.ram_block1a20(\ram_block1a20~PORTBDATAOUT0 ),
	.ram_block1a85(\ram_block1a85~PORTBDATAOUT0 ),
	.ram_block1a21(\ram_block1a21~PORTBDATAOUT0 ),
	.ram_block1a86(\ram_block1a86~PORTBDATAOUT0 ),
	.ram_block1a22(\ram_block1a22~PORTBDATAOUT0 ),
	.ram_block1a87(\ram_block1a87~PORTBDATAOUT0 ),
	.ram_block1a23(\ram_block1a23~PORTBDATAOUT0 ),
	.ram_block1a88(\ram_block1a88~PORTBDATAOUT0 ),
	.ram_block1a24(\ram_block1a24~PORTBDATAOUT0 ),
	.ram_block1a89(\ram_block1a89~PORTBDATAOUT0 ),
	.ram_block1a25(\ram_block1a25~PORTBDATAOUT0 ),
	.ram_block1a90(\ram_block1a90~PORTBDATAOUT0 ),
	.ram_block1a26(\ram_block1a26~PORTBDATAOUT0 ),
	.ram_block1a91(\ram_block1a91~PORTBDATAOUT0 ),
	.ram_block1a27(\ram_block1a27~PORTBDATAOUT0 ),
	.ram_block1a92(\ram_block1a92~PORTBDATAOUT0 ),
	.ram_block1a28(\ram_block1a28~PORTBDATAOUT0 ),
	.ram_block1a93(\ram_block1a93~PORTBDATAOUT0 ),
	.ram_block1a29(\ram_block1a29~PORTBDATAOUT0 ),
	.ram_block1a94(\ram_block1a94~PORTBDATAOUT0 ),
	.ram_block1a30(\ram_block1a30~PORTBDATAOUT0 ),
	.ram_block1a95(\ram_block1a95~PORTBDATAOUT0 ),
	.ram_block1a31(\ram_block1a31~PORTBDATAOUT0 ),
	.ram_block1a96(\ram_block1a96~PORTBDATAOUT0 ),
	.ram_block1a32(\ram_block1a32~PORTBDATAOUT0 ),
	.ram_block1a97(\ram_block1a97~PORTBDATAOUT0 ),
	.ram_block1a33(\ram_block1a33~PORTBDATAOUT0 ),
	.ram_block1a98(\ram_block1a98~PORTBDATAOUT0 ),
	.ram_block1a34(\ram_block1a34~PORTBDATAOUT0 ),
	.ram_block1a99(\ram_block1a99~PORTBDATAOUT0 ),
	.ram_block1a35(\ram_block1a35~PORTBDATAOUT0 ),
	.ram_block1a100(\ram_block1a100~PORTBDATAOUT0 ),
	.ram_block1a36(\ram_block1a36~PORTBDATAOUT0 ),
	.ram_block1a101(\ram_block1a101~PORTBDATAOUT0 ),
	.ram_block1a37(\ram_block1a37~PORTBDATAOUT0 ),
	.ram_block1a102(\ram_block1a102~PORTBDATAOUT0 ),
	.ram_block1a38(\ram_block1a38~PORTBDATAOUT0 ),
	.ram_block1a103(\ram_block1a103~PORTBDATAOUT0 ),
	.ram_block1a39(\ram_block1a39~PORTBDATAOUT0 ),
	.ram_block1a104(\ram_block1a104~PORTBDATAOUT0 ),
	.ram_block1a40(\ram_block1a40~PORTBDATAOUT0 ),
	.ram_block1a105(\ram_block1a105~PORTBDATAOUT0 ),
	.ram_block1a41(\ram_block1a41~PORTBDATAOUT0 ),
	.ram_block1a106(\ram_block1a106~PORTBDATAOUT0 ),
	.ram_block1a42(\ram_block1a42~PORTBDATAOUT0 ),
	.ram_block1a107(\ram_block1a107~PORTBDATAOUT0 ),
	.ram_block1a43(\ram_block1a43~PORTBDATAOUT0 ),
	.ram_block1a108(\ram_block1a108~PORTBDATAOUT0 ),
	.ram_block1a44(\ram_block1a44~PORTBDATAOUT0 ),
	.ram_block1a109(\ram_block1a109~PORTBDATAOUT0 ),
	.ram_block1a45(\ram_block1a45~PORTBDATAOUT0 ),
	.ram_block1a110(\ram_block1a110~PORTBDATAOUT0 ),
	.ram_block1a46(\ram_block1a46~PORTBDATAOUT0 ),
	.ram_block1a111(\ram_block1a111~PORTBDATAOUT0 ),
	.ram_block1a47(\ram_block1a47~PORTBDATAOUT0 ),
	.ram_block1a112(\ram_block1a112~PORTBDATAOUT0 ),
	.ram_block1a48(\ram_block1a48~PORTBDATAOUT0 ),
	.ram_block1a113(\ram_block1a113~PORTBDATAOUT0 ),
	.ram_block1a49(\ram_block1a49~PORTBDATAOUT0 ),
	.ram_block1a114(\ram_block1a114~PORTBDATAOUT0 ),
	.ram_block1a50(\ram_block1a50~PORTBDATAOUT0 ),
	.ram_block1a115(\ram_block1a115~PORTBDATAOUT0 ),
	.ram_block1a51(\ram_block1a51~PORTBDATAOUT0 ),
	.ram_block1a116(\ram_block1a116~PORTBDATAOUT0 ),
	.ram_block1a52(\ram_block1a52~PORTBDATAOUT0 ),
	.ram_block1a117(\ram_block1a117~PORTBDATAOUT0 ),
	.ram_block1a53(\ram_block1a53~PORTBDATAOUT0 ),
	.ram_block1a118(\ram_block1a118~PORTBDATAOUT0 ),
	.ram_block1a54(\ram_block1a54~PORTBDATAOUT0 ),
	.ram_block1a119(\ram_block1a119~PORTBDATAOUT0 ),
	.ram_block1a55(\ram_block1a55~PORTBDATAOUT0 ),
	.ram_block1a120(\ram_block1a120~PORTBDATAOUT0 ),
	.ram_block1a56(\ram_block1a56~PORTBDATAOUT0 ),
	.ram_block1a121(\ram_block1a121~PORTBDATAOUT0 ),
	.ram_block1a57(\ram_block1a57~PORTBDATAOUT0 ),
	.ram_block1a122(\ram_block1a122~PORTBDATAOUT0 ),
	.ram_block1a58(\ram_block1a58~PORTBDATAOUT0 ),
	.ram_block1a123(\ram_block1a123~PORTBDATAOUT0 ),
	.ram_block1a59(\ram_block1a59~PORTBDATAOUT0 ),
	.ram_block1a124(\ram_block1a124~PORTBDATAOUT0 ),
	.ram_block1a60(\ram_block1a60~PORTBDATAOUT0 ),
	.ram_block1a125(\ram_block1a125~PORTBDATAOUT0 ),
	.ram_block1a61(\ram_block1a61~PORTBDATAOUT0 ),
	.ram_block1a126(\ram_block1a126~PORTBDATAOUT0 ),
	.ram_block1a62(\ram_block1a62~PORTBDATAOUT0 ),
	.ram_block1a127(\ram_block1a127~PORTBDATAOUT0 ),
	.ram_block1a63(\ram_block1a63~PORTBDATAOUT0 ),
	.address_reg_b_0(\address_reg_b[0]~q ),
	.result_node_0(result_node_01),
	.result_node_1(result_node_110),
	.result_node_2(result_node_210),
	.result_node_3(result_node_310),
	.result_node_4(result_node_410),
	.result_node_5(result_node_510),
	.result_node_6(result_node_64),
	.result_node_7(result_node_71),
	.result_node_8(result_node_81),
	.result_node_9(result_node_91),
	.result_node_10(result_node_101),
	.result_node_11(result_node_111),
	.result_node_12(result_node_121),
	.result_node_13(result_node_131),
	.result_node_14(result_node_141),
	.result_node_15(result_node_151),
	.result_node_16(result_node_161),
	.result_node_17(result_node_171),
	.result_node_18(result_node_181),
	.result_node_19(result_node_191),
	.result_node_20(result_node_201),
	.result_node_21(result_node_211),
	.result_node_22(result_node_221),
	.result_node_23(result_node_231),
	.result_node_24(result_node_241),
	.result_node_25(result_node_251),
	.result_node_26(result_node_261),
	.result_node_27(result_node_271),
	.result_node_28(result_node_281),
	.result_node_29(result_node_291),
	.result_node_30(result_node_301),
	.result_node_31(result_node_311),
	.result_node_32(result_node_321),
	.result_node_33(result_node_331),
	.result_node_34(result_node_341),
	.result_node_35(result_node_351),
	.result_node_36(result_node_361),
	.result_node_37(result_node_371),
	.result_node_38(result_node_381),
	.result_node_39(result_node_391),
	.result_node_40(result_node_401),
	.result_node_41(result_node_411),
	.result_node_42(result_node_421),
	.result_node_43(result_node_431),
	.result_node_44(result_node_441),
	.result_node_45(result_node_451),
	.result_node_46(result_node_461),
	.result_node_47(result_node_471),
	.result_node_48(result_node_481),
	.result_node_49(result_node_491),
	.result_node_50(result_node_501),
	.result_node_51(result_node_511),
	.result_node_52(result_node_521),
	.result_node_53(result_node_531),
	.result_node_54(result_node_541),
	.result_node_55(result_node_551),
	.result_node_56(result_node_561),
	.result_node_57(result_node_571),
	.result_node_58(result_node_581),
	.result_node_59(result_node_591),
	.result_node_60(result_node_601),
	.result_node_61(result_node_611),
	.result_node_62(result_node_621),
	.result_node_63(result_node_631));

qtestpd_mux_fsb mux4(
	.ram_block1a64(\ram_block1a64~portadataout ),
	.ram_block1a0(\ram_block1a0~portadataout ),
	.ram_block1a65(\ram_block1a65~portadataout ),
	.ram_block1a1(\ram_block1a1~portadataout ),
	.ram_block1a66(\ram_block1a66~portadataout ),
	.ram_block1a2(\ram_block1a2~portadataout ),
	.ram_block1a67(\ram_block1a67~portadataout ),
	.ram_block1a3(\ram_block1a3~portadataout ),
	.ram_block1a68(\ram_block1a68~portadataout ),
	.ram_block1a4(\ram_block1a4~portadataout ),
	.ram_block1a69(\ram_block1a69~portadataout ),
	.ram_block1a5(\ram_block1a5~portadataout ),
	.ram_block1a70(\ram_block1a70~portadataout ),
	.ram_block1a6(\ram_block1a6~portadataout ),
	.ram_block1a71(\ram_block1a71~portadataout ),
	.ram_block1a7(\ram_block1a7~portadataout ),
	.ram_block1a72(\ram_block1a72~portadataout ),
	.ram_block1a8(\ram_block1a8~portadataout ),
	.ram_block1a73(\ram_block1a73~portadataout ),
	.ram_block1a9(\ram_block1a9~portadataout ),
	.ram_block1a74(\ram_block1a74~portadataout ),
	.ram_block1a10(\ram_block1a10~portadataout ),
	.ram_block1a75(\ram_block1a75~portadataout ),
	.ram_block1a11(\ram_block1a11~portadataout ),
	.ram_block1a76(\ram_block1a76~portadataout ),
	.ram_block1a12(\ram_block1a12~portadataout ),
	.ram_block1a77(\ram_block1a77~portadataout ),
	.ram_block1a13(\ram_block1a13~portadataout ),
	.ram_block1a78(\ram_block1a78~portadataout ),
	.ram_block1a14(\ram_block1a14~portadataout ),
	.ram_block1a79(\ram_block1a79~portadataout ),
	.ram_block1a15(\ram_block1a15~portadataout ),
	.ram_block1a80(\ram_block1a80~portadataout ),
	.ram_block1a16(\ram_block1a16~portadataout ),
	.ram_block1a81(\ram_block1a81~portadataout ),
	.ram_block1a17(\ram_block1a17~portadataout ),
	.ram_block1a82(\ram_block1a82~portadataout ),
	.ram_block1a18(\ram_block1a18~portadataout ),
	.ram_block1a83(\ram_block1a83~portadataout ),
	.ram_block1a19(\ram_block1a19~portadataout ),
	.ram_block1a84(\ram_block1a84~portadataout ),
	.ram_block1a20(\ram_block1a20~portadataout ),
	.ram_block1a85(\ram_block1a85~portadataout ),
	.ram_block1a21(\ram_block1a21~portadataout ),
	.ram_block1a86(\ram_block1a86~portadataout ),
	.ram_block1a22(\ram_block1a22~portadataout ),
	.ram_block1a87(\ram_block1a87~portadataout ),
	.ram_block1a23(\ram_block1a23~portadataout ),
	.ram_block1a88(\ram_block1a88~portadataout ),
	.ram_block1a24(\ram_block1a24~portadataout ),
	.ram_block1a89(\ram_block1a89~portadataout ),
	.ram_block1a25(\ram_block1a25~portadataout ),
	.ram_block1a90(\ram_block1a90~portadataout ),
	.ram_block1a26(\ram_block1a26~portadataout ),
	.ram_block1a91(\ram_block1a91~portadataout ),
	.ram_block1a27(\ram_block1a27~portadataout ),
	.ram_block1a92(\ram_block1a92~portadataout ),
	.ram_block1a28(\ram_block1a28~portadataout ),
	.ram_block1a93(\ram_block1a93~portadataout ),
	.ram_block1a29(\ram_block1a29~portadataout ),
	.ram_block1a94(\ram_block1a94~portadataout ),
	.ram_block1a30(\ram_block1a30~portadataout ),
	.ram_block1a95(\ram_block1a95~portadataout ),
	.ram_block1a31(\ram_block1a31~portadataout ),
	.ram_block1a96(\ram_block1a96~portadataout ),
	.ram_block1a32(\ram_block1a32~portadataout ),
	.ram_block1a97(\ram_block1a97~portadataout ),
	.ram_block1a33(\ram_block1a33~portadataout ),
	.ram_block1a98(\ram_block1a98~portadataout ),
	.ram_block1a34(\ram_block1a34~portadataout ),
	.ram_block1a99(\ram_block1a99~portadataout ),
	.ram_block1a35(\ram_block1a35~portadataout ),
	.ram_block1a100(\ram_block1a100~portadataout ),
	.ram_block1a36(\ram_block1a36~portadataout ),
	.ram_block1a101(\ram_block1a101~portadataout ),
	.ram_block1a37(\ram_block1a37~portadataout ),
	.ram_block1a102(\ram_block1a102~portadataout ),
	.ram_block1a38(\ram_block1a38~portadataout ),
	.ram_block1a103(\ram_block1a103~portadataout ),
	.ram_block1a39(\ram_block1a39~portadataout ),
	.ram_block1a104(\ram_block1a104~portadataout ),
	.ram_block1a40(\ram_block1a40~portadataout ),
	.ram_block1a105(\ram_block1a105~portadataout ),
	.ram_block1a41(\ram_block1a41~portadataout ),
	.ram_block1a106(\ram_block1a106~portadataout ),
	.ram_block1a42(\ram_block1a42~portadataout ),
	.ram_block1a107(\ram_block1a107~portadataout ),
	.ram_block1a43(\ram_block1a43~portadataout ),
	.ram_block1a108(\ram_block1a108~portadataout ),
	.ram_block1a44(\ram_block1a44~portadataout ),
	.ram_block1a109(\ram_block1a109~portadataout ),
	.ram_block1a45(\ram_block1a45~portadataout ),
	.ram_block1a110(\ram_block1a110~portadataout ),
	.ram_block1a46(\ram_block1a46~portadataout ),
	.ram_block1a111(\ram_block1a111~portadataout ),
	.ram_block1a47(\ram_block1a47~portadataout ),
	.ram_block1a112(\ram_block1a112~portadataout ),
	.ram_block1a48(\ram_block1a48~portadataout ),
	.ram_block1a113(\ram_block1a113~portadataout ),
	.ram_block1a49(\ram_block1a49~portadataout ),
	.ram_block1a114(\ram_block1a114~portadataout ),
	.ram_block1a50(\ram_block1a50~portadataout ),
	.ram_block1a115(\ram_block1a115~portadataout ),
	.ram_block1a51(\ram_block1a51~portadataout ),
	.ram_block1a116(\ram_block1a116~portadataout ),
	.ram_block1a52(\ram_block1a52~portadataout ),
	.ram_block1a117(\ram_block1a117~portadataout ),
	.ram_block1a53(\ram_block1a53~portadataout ),
	.ram_block1a118(\ram_block1a118~portadataout ),
	.ram_block1a54(\ram_block1a54~portadataout ),
	.ram_block1a119(\ram_block1a119~portadataout ),
	.ram_block1a55(\ram_block1a55~portadataout ),
	.ram_block1a120(\ram_block1a120~portadataout ),
	.ram_block1a56(\ram_block1a56~portadataout ),
	.ram_block1a121(\ram_block1a121~portadataout ),
	.ram_block1a57(\ram_block1a57~portadataout ),
	.ram_block1a122(\ram_block1a122~portadataout ),
	.ram_block1a58(\ram_block1a58~portadataout ),
	.ram_block1a123(\ram_block1a123~portadataout ),
	.ram_block1a59(\ram_block1a59~portadataout ),
	.ram_block1a124(\ram_block1a124~portadataout ),
	.ram_block1a60(\ram_block1a60~portadataout ),
	.ram_block1a125(\ram_block1a125~portadataout ),
	.ram_block1a61(\ram_block1a61~portadataout ),
	.ram_block1a126(\ram_block1a126~portadataout ),
	.ram_block1a62(\ram_block1a62~portadataout ),
	.ram_block1a127(\ram_block1a127~portadataout ),
	.ram_block1a63(\ram_block1a63~portadataout ),
	.address_reg_a_0(\address_reg_a[0]~q ),
	.result_node_0(result_node_0),
	.result_node_1(result_node_1),
	.result_node_2(result_node_2),
	.result_node_3(result_node_3),
	.result_node_4(result_node_4),
	.result_node_5(result_node_5),
	.result_node_6(result_node_6),
	.result_node_7(result_node_7),
	.result_node_8(result_node_8),
	.result_node_9(result_node_9),
	.result_node_10(result_node_10),
	.result_node_11(result_node_11),
	.result_node_12(result_node_12),
	.result_node_13(result_node_13),
	.result_node_14(result_node_14),
	.result_node_15(result_node_15),
	.result_node_16(result_node_16),
	.result_node_17(result_node_17),
	.result_node_18(result_node_18),
	.result_node_19(result_node_19),
	.result_node_20(result_node_20),
	.result_node_21(result_node_21),
	.result_node_22(result_node_22),
	.result_node_23(result_node_23),
	.result_node_24(result_node_24),
	.result_node_25(result_node_25),
	.result_node_26(result_node_26),
	.result_node_27(result_node_27),
	.result_node_28(result_node_28),
	.result_node_29(result_node_29),
	.result_node_30(result_node_30),
	.result_node_31(result_node_31),
	.result_node_32(result_node_32),
	.result_node_33(result_node_33),
	.result_node_34(result_node_34),
	.result_node_35(result_node_35),
	.result_node_36(result_node_36),
	.result_node_37(result_node_37),
	.result_node_38(result_node_38),
	.result_node_39(result_node_39),
	.result_node_40(result_node_40),
	.result_node_41(result_node_41),
	.result_node_42(result_node_42),
	.result_node_43(result_node_43),
	.result_node_44(result_node_44),
	.result_node_45(result_node_45),
	.result_node_46(result_node_46),
	.result_node_47(result_node_47),
	.result_node_48(result_node_48),
	.result_node_49(result_node_49),
	.result_node_50(result_node_50),
	.result_node_51(result_node_51),
	.result_node_52(result_node_52),
	.result_node_53(result_node_53),
	.result_node_54(result_node_54),
	.result_node_55(result_node_55),
	.result_node_56(result_node_56),
	.result_node_57(result_node_57),
	.result_node_58(result_node_58),
	.result_node_59(result_node_59),
	.result_node_60(result_node_60),
	.result_node_61(result_node_61),
	.result_node_62(result_node_62),
	.result_node_63(result_node_63));

qtestpd_decode_d0b_1 decode3(
	.eq_node_1(\decode3|eq_node[1]~0_combout ),
	.eq_node_0(\decode3|eq_node[0]~1_combout ),
	.onchip_memory2_0_s2_address_13(address_b[13]),
	.onchip_memory2_0_s2_chipselect(onchip_memory2_0_s2_chipselect),
	.onchip_memory2_0_s2_write(onchip_memory2_0_s2_write));

qtestpd_decode_d0b decode2(
	.eq_node_1(\decode2|eq_node[1]~0_combout ),
	.eq_node_0(\decode2|eq_node[0]~1_combout ),
	.onchip_memory2_0_s1_address_13(address_a[13]),
	.onchip_memory2_0_s1_chipselect(onchip_memory2_0_s1_chipselect),
	.onchip_memory2_0_s1_write(onchip_memory2_0_s1_write));

cycloneiv_ram_block ram_block1a64(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[0]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a64_PORTADATAOUT_bus),
	.portbdataout(ram_block1a64_PORTBDATAOUT_bus));
defparam ram_block1a64.clk0_core_clock_enable = "ena0";
defparam ram_block1a64.clk0_input_clock_enable = "ena0";
defparam ram_block1a64.clk1_core_clock_enable = "ena1";
defparam ram_block1a64.clk1_input_clock_enable = "ena1";
defparam ram_block1a64.data_interleave_offset_in_bits = 1;
defparam ram_block1a64.data_interleave_width_in_bits = 1;
defparam ram_block1a64.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a64.init_file_layout = "port_a";
defparam ram_block1a64.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a64.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a64.operation_mode = "bidir_dual_port";
defparam ram_block1a64.port_a_address_clear = "none";
defparam ram_block1a64.port_a_address_width = 13;
defparam ram_block1a64.port_a_byte_enable_mask_width = 1;
defparam ram_block1a64.port_a_byte_size = 1;
defparam ram_block1a64.port_a_data_out_clear = "none";
defparam ram_block1a64.port_a_data_out_clock = "none";
defparam ram_block1a64.port_a_data_width = 1;
defparam ram_block1a64.port_a_first_address = 8192;
defparam ram_block1a64.port_a_first_bit_number = 0;
defparam ram_block1a64.port_a_last_address = 16383;
defparam ram_block1a64.port_a_logical_ram_depth = 16384;
defparam ram_block1a64.port_a_logical_ram_width = 64;
defparam ram_block1a64.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a64.port_b_address_clear = "none";
defparam ram_block1a64.port_b_address_clock = "clock1";
defparam ram_block1a64.port_b_address_width = 13;
defparam ram_block1a64.port_b_byte_enable_clock = "clock1";
defparam ram_block1a64.port_b_byte_enable_mask_width = 1;
defparam ram_block1a64.port_b_byte_size = 1;
defparam ram_block1a64.port_b_data_in_clock = "clock1";
defparam ram_block1a64.port_b_data_out_clear = "none";
defparam ram_block1a64.port_b_data_out_clock = "none";
defparam ram_block1a64.port_b_data_width = 1;
defparam ram_block1a64.port_b_first_address = 8192;
defparam ram_block1a64.port_b_first_bit_number = 0;
defparam ram_block1a64.port_b_last_address = 16383;
defparam ram_block1a64.port_b_logical_ram_depth = 16384;
defparam ram_block1a64.port_b_logical_ram_width = 64;
defparam ram_block1a64.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a64.port_b_read_enable_clock = "clock1";
defparam ram_block1a64.port_b_write_enable_clock = "clock1";
defparam ram_block1a64.ram_block_type = "auto";
defparam ram_block1a64.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a64.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a64.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a64.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a0(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[0]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.clk1_input_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "bidir_dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 13;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 8191;
defparam ram_block1a0.port_a_logical_ram_depth = 16384;
defparam ram_block1a0.port_a_logical_ram_width = 64;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 13;
defparam ram_block1a0.port_b_byte_enable_clock = "clock1";
defparam ram_block1a0.port_b_byte_enable_mask_width = 1;
defparam ram_block1a0.port_b_byte_size = 1;
defparam ram_block1a0.port_b_data_in_clock = "clock1";
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 8191;
defparam ram_block1a0.port_b_logical_ram_depth = 16384;
defparam ram_block1a0.port_b_logical_ram_width = 64;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.port_b_write_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a0.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a65(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[1]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a65_PORTADATAOUT_bus),
	.portbdataout(ram_block1a65_PORTBDATAOUT_bus));
defparam ram_block1a65.clk0_core_clock_enable = "ena0";
defparam ram_block1a65.clk0_input_clock_enable = "ena0";
defparam ram_block1a65.clk1_core_clock_enable = "ena1";
defparam ram_block1a65.clk1_input_clock_enable = "ena1";
defparam ram_block1a65.data_interleave_offset_in_bits = 1;
defparam ram_block1a65.data_interleave_width_in_bits = 1;
defparam ram_block1a65.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a65.init_file_layout = "port_a";
defparam ram_block1a65.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a65.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a65.operation_mode = "bidir_dual_port";
defparam ram_block1a65.port_a_address_clear = "none";
defparam ram_block1a65.port_a_address_width = 13;
defparam ram_block1a65.port_a_byte_enable_mask_width = 1;
defparam ram_block1a65.port_a_byte_size = 1;
defparam ram_block1a65.port_a_data_out_clear = "none";
defparam ram_block1a65.port_a_data_out_clock = "none";
defparam ram_block1a65.port_a_data_width = 1;
defparam ram_block1a65.port_a_first_address = 8192;
defparam ram_block1a65.port_a_first_bit_number = 1;
defparam ram_block1a65.port_a_last_address = 16383;
defparam ram_block1a65.port_a_logical_ram_depth = 16384;
defparam ram_block1a65.port_a_logical_ram_width = 64;
defparam ram_block1a65.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a65.port_b_address_clear = "none";
defparam ram_block1a65.port_b_address_clock = "clock1";
defparam ram_block1a65.port_b_address_width = 13;
defparam ram_block1a65.port_b_byte_enable_clock = "clock1";
defparam ram_block1a65.port_b_byte_enable_mask_width = 1;
defparam ram_block1a65.port_b_byte_size = 1;
defparam ram_block1a65.port_b_data_in_clock = "clock1";
defparam ram_block1a65.port_b_data_out_clear = "none";
defparam ram_block1a65.port_b_data_out_clock = "none";
defparam ram_block1a65.port_b_data_width = 1;
defparam ram_block1a65.port_b_first_address = 8192;
defparam ram_block1a65.port_b_first_bit_number = 1;
defparam ram_block1a65.port_b_last_address = 16383;
defparam ram_block1a65.port_b_logical_ram_depth = 16384;
defparam ram_block1a65.port_b_logical_ram_width = 64;
defparam ram_block1a65.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a65.port_b_read_enable_clock = "clock1";
defparam ram_block1a65.port_b_write_enable_clock = "clock1";
defparam ram_block1a65.ram_block_type = "auto";
defparam ram_block1a65.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a65.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a65.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a65.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a1(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[1]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.clk1_input_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "bidir_dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 13;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 8191;
defparam ram_block1a1.port_a_logical_ram_depth = 16384;
defparam ram_block1a1.port_a_logical_ram_width = 64;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 13;
defparam ram_block1a1.port_b_byte_enable_clock = "clock1";
defparam ram_block1a1.port_b_byte_enable_mask_width = 1;
defparam ram_block1a1.port_b_byte_size = 1;
defparam ram_block1a1.port_b_data_in_clock = "clock1";
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 8191;
defparam ram_block1a1.port_b_logical_ram_depth = 16384;
defparam ram_block1a1.port_b_logical_ram_width = 64;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.port_b_write_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a1.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a66(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[2]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a66_PORTADATAOUT_bus),
	.portbdataout(ram_block1a66_PORTBDATAOUT_bus));
defparam ram_block1a66.clk0_core_clock_enable = "ena0";
defparam ram_block1a66.clk0_input_clock_enable = "ena0";
defparam ram_block1a66.clk1_core_clock_enable = "ena1";
defparam ram_block1a66.clk1_input_clock_enable = "ena1";
defparam ram_block1a66.data_interleave_offset_in_bits = 1;
defparam ram_block1a66.data_interleave_width_in_bits = 1;
defparam ram_block1a66.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a66.init_file_layout = "port_a";
defparam ram_block1a66.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a66.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a66.operation_mode = "bidir_dual_port";
defparam ram_block1a66.port_a_address_clear = "none";
defparam ram_block1a66.port_a_address_width = 13;
defparam ram_block1a66.port_a_byte_enable_mask_width = 1;
defparam ram_block1a66.port_a_byte_size = 1;
defparam ram_block1a66.port_a_data_out_clear = "none";
defparam ram_block1a66.port_a_data_out_clock = "none";
defparam ram_block1a66.port_a_data_width = 1;
defparam ram_block1a66.port_a_first_address = 8192;
defparam ram_block1a66.port_a_first_bit_number = 2;
defparam ram_block1a66.port_a_last_address = 16383;
defparam ram_block1a66.port_a_logical_ram_depth = 16384;
defparam ram_block1a66.port_a_logical_ram_width = 64;
defparam ram_block1a66.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a66.port_b_address_clear = "none";
defparam ram_block1a66.port_b_address_clock = "clock1";
defparam ram_block1a66.port_b_address_width = 13;
defparam ram_block1a66.port_b_byte_enable_clock = "clock1";
defparam ram_block1a66.port_b_byte_enable_mask_width = 1;
defparam ram_block1a66.port_b_byte_size = 1;
defparam ram_block1a66.port_b_data_in_clock = "clock1";
defparam ram_block1a66.port_b_data_out_clear = "none";
defparam ram_block1a66.port_b_data_out_clock = "none";
defparam ram_block1a66.port_b_data_width = 1;
defparam ram_block1a66.port_b_first_address = 8192;
defparam ram_block1a66.port_b_first_bit_number = 2;
defparam ram_block1a66.port_b_last_address = 16383;
defparam ram_block1a66.port_b_logical_ram_depth = 16384;
defparam ram_block1a66.port_b_logical_ram_width = 64;
defparam ram_block1a66.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a66.port_b_read_enable_clock = "clock1";
defparam ram_block1a66.port_b_write_enable_clock = "clock1";
defparam ram_block1a66.ram_block_type = "auto";
defparam ram_block1a66.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a66.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a66.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a66.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a2(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[2]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.clk1_input_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "bidir_dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 13;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 8191;
defparam ram_block1a2.port_a_logical_ram_depth = 16384;
defparam ram_block1a2.port_a_logical_ram_width = 64;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 13;
defparam ram_block1a2.port_b_byte_enable_clock = "clock1";
defparam ram_block1a2.port_b_byte_enable_mask_width = 1;
defparam ram_block1a2.port_b_byte_size = 1;
defparam ram_block1a2.port_b_data_in_clock = "clock1";
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 8191;
defparam ram_block1a2.port_b_logical_ram_depth = 16384;
defparam ram_block1a2.port_b_logical_ram_width = 64;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.port_b_write_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a2.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a67(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[3]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a67_PORTADATAOUT_bus),
	.portbdataout(ram_block1a67_PORTBDATAOUT_bus));
defparam ram_block1a67.clk0_core_clock_enable = "ena0";
defparam ram_block1a67.clk0_input_clock_enable = "ena0";
defparam ram_block1a67.clk1_core_clock_enable = "ena1";
defparam ram_block1a67.clk1_input_clock_enable = "ena1";
defparam ram_block1a67.data_interleave_offset_in_bits = 1;
defparam ram_block1a67.data_interleave_width_in_bits = 1;
defparam ram_block1a67.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a67.init_file_layout = "port_a";
defparam ram_block1a67.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a67.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a67.operation_mode = "bidir_dual_port";
defparam ram_block1a67.port_a_address_clear = "none";
defparam ram_block1a67.port_a_address_width = 13;
defparam ram_block1a67.port_a_byte_enable_mask_width = 1;
defparam ram_block1a67.port_a_byte_size = 1;
defparam ram_block1a67.port_a_data_out_clear = "none";
defparam ram_block1a67.port_a_data_out_clock = "none";
defparam ram_block1a67.port_a_data_width = 1;
defparam ram_block1a67.port_a_first_address = 8192;
defparam ram_block1a67.port_a_first_bit_number = 3;
defparam ram_block1a67.port_a_last_address = 16383;
defparam ram_block1a67.port_a_logical_ram_depth = 16384;
defparam ram_block1a67.port_a_logical_ram_width = 64;
defparam ram_block1a67.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a67.port_b_address_clear = "none";
defparam ram_block1a67.port_b_address_clock = "clock1";
defparam ram_block1a67.port_b_address_width = 13;
defparam ram_block1a67.port_b_byte_enable_clock = "clock1";
defparam ram_block1a67.port_b_byte_enable_mask_width = 1;
defparam ram_block1a67.port_b_byte_size = 1;
defparam ram_block1a67.port_b_data_in_clock = "clock1";
defparam ram_block1a67.port_b_data_out_clear = "none";
defparam ram_block1a67.port_b_data_out_clock = "none";
defparam ram_block1a67.port_b_data_width = 1;
defparam ram_block1a67.port_b_first_address = 8192;
defparam ram_block1a67.port_b_first_bit_number = 3;
defparam ram_block1a67.port_b_last_address = 16383;
defparam ram_block1a67.port_b_logical_ram_depth = 16384;
defparam ram_block1a67.port_b_logical_ram_width = 64;
defparam ram_block1a67.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a67.port_b_read_enable_clock = "clock1";
defparam ram_block1a67.port_b_write_enable_clock = "clock1";
defparam ram_block1a67.ram_block_type = "auto";
defparam ram_block1a67.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a67.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a67.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a67.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a3(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[3]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.clk1_input_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "bidir_dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 13;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 8191;
defparam ram_block1a3.port_a_logical_ram_depth = 16384;
defparam ram_block1a3.port_a_logical_ram_width = 64;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 13;
defparam ram_block1a3.port_b_byte_enable_clock = "clock1";
defparam ram_block1a3.port_b_byte_enable_mask_width = 1;
defparam ram_block1a3.port_b_byte_size = 1;
defparam ram_block1a3.port_b_data_in_clock = "clock1";
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 8191;
defparam ram_block1a3.port_b_logical_ram_depth = 16384;
defparam ram_block1a3.port_b_logical_ram_width = 64;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.port_b_write_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a3.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a68(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[4]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a68_PORTADATAOUT_bus),
	.portbdataout(ram_block1a68_PORTBDATAOUT_bus));
defparam ram_block1a68.clk0_core_clock_enable = "ena0";
defparam ram_block1a68.clk0_input_clock_enable = "ena0";
defparam ram_block1a68.clk1_core_clock_enable = "ena1";
defparam ram_block1a68.clk1_input_clock_enable = "ena1";
defparam ram_block1a68.data_interleave_offset_in_bits = 1;
defparam ram_block1a68.data_interleave_width_in_bits = 1;
defparam ram_block1a68.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a68.init_file_layout = "port_a";
defparam ram_block1a68.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a68.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a68.operation_mode = "bidir_dual_port";
defparam ram_block1a68.port_a_address_clear = "none";
defparam ram_block1a68.port_a_address_width = 13;
defparam ram_block1a68.port_a_byte_enable_mask_width = 1;
defparam ram_block1a68.port_a_byte_size = 1;
defparam ram_block1a68.port_a_data_out_clear = "none";
defparam ram_block1a68.port_a_data_out_clock = "none";
defparam ram_block1a68.port_a_data_width = 1;
defparam ram_block1a68.port_a_first_address = 8192;
defparam ram_block1a68.port_a_first_bit_number = 4;
defparam ram_block1a68.port_a_last_address = 16383;
defparam ram_block1a68.port_a_logical_ram_depth = 16384;
defparam ram_block1a68.port_a_logical_ram_width = 64;
defparam ram_block1a68.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a68.port_b_address_clear = "none";
defparam ram_block1a68.port_b_address_clock = "clock1";
defparam ram_block1a68.port_b_address_width = 13;
defparam ram_block1a68.port_b_byte_enable_clock = "clock1";
defparam ram_block1a68.port_b_byte_enable_mask_width = 1;
defparam ram_block1a68.port_b_byte_size = 1;
defparam ram_block1a68.port_b_data_in_clock = "clock1";
defparam ram_block1a68.port_b_data_out_clear = "none";
defparam ram_block1a68.port_b_data_out_clock = "none";
defparam ram_block1a68.port_b_data_width = 1;
defparam ram_block1a68.port_b_first_address = 8192;
defparam ram_block1a68.port_b_first_bit_number = 4;
defparam ram_block1a68.port_b_last_address = 16383;
defparam ram_block1a68.port_b_logical_ram_depth = 16384;
defparam ram_block1a68.port_b_logical_ram_width = 64;
defparam ram_block1a68.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a68.port_b_read_enable_clock = "clock1";
defparam ram_block1a68.port_b_write_enable_clock = "clock1";
defparam ram_block1a68.ram_block_type = "auto";
defparam ram_block1a68.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a68.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a68.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a68.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a4(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[4]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.clk1_input_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "bidir_dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 13;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 8191;
defparam ram_block1a4.port_a_logical_ram_depth = 16384;
defparam ram_block1a4.port_a_logical_ram_width = 64;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 13;
defparam ram_block1a4.port_b_byte_enable_clock = "clock1";
defparam ram_block1a4.port_b_byte_enable_mask_width = 1;
defparam ram_block1a4.port_b_byte_size = 1;
defparam ram_block1a4.port_b_data_in_clock = "clock1";
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 8191;
defparam ram_block1a4.port_b_logical_ram_depth = 16384;
defparam ram_block1a4.port_b_logical_ram_width = 64;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.port_b_write_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a4.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a69(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[5]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a69_PORTADATAOUT_bus),
	.portbdataout(ram_block1a69_PORTBDATAOUT_bus));
defparam ram_block1a69.clk0_core_clock_enable = "ena0";
defparam ram_block1a69.clk0_input_clock_enable = "ena0";
defparam ram_block1a69.clk1_core_clock_enable = "ena1";
defparam ram_block1a69.clk1_input_clock_enable = "ena1";
defparam ram_block1a69.data_interleave_offset_in_bits = 1;
defparam ram_block1a69.data_interleave_width_in_bits = 1;
defparam ram_block1a69.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a69.init_file_layout = "port_a";
defparam ram_block1a69.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a69.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a69.operation_mode = "bidir_dual_port";
defparam ram_block1a69.port_a_address_clear = "none";
defparam ram_block1a69.port_a_address_width = 13;
defparam ram_block1a69.port_a_byte_enable_mask_width = 1;
defparam ram_block1a69.port_a_byte_size = 1;
defparam ram_block1a69.port_a_data_out_clear = "none";
defparam ram_block1a69.port_a_data_out_clock = "none";
defparam ram_block1a69.port_a_data_width = 1;
defparam ram_block1a69.port_a_first_address = 8192;
defparam ram_block1a69.port_a_first_bit_number = 5;
defparam ram_block1a69.port_a_last_address = 16383;
defparam ram_block1a69.port_a_logical_ram_depth = 16384;
defparam ram_block1a69.port_a_logical_ram_width = 64;
defparam ram_block1a69.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a69.port_b_address_clear = "none";
defparam ram_block1a69.port_b_address_clock = "clock1";
defparam ram_block1a69.port_b_address_width = 13;
defparam ram_block1a69.port_b_byte_enable_clock = "clock1";
defparam ram_block1a69.port_b_byte_enable_mask_width = 1;
defparam ram_block1a69.port_b_byte_size = 1;
defparam ram_block1a69.port_b_data_in_clock = "clock1";
defparam ram_block1a69.port_b_data_out_clear = "none";
defparam ram_block1a69.port_b_data_out_clock = "none";
defparam ram_block1a69.port_b_data_width = 1;
defparam ram_block1a69.port_b_first_address = 8192;
defparam ram_block1a69.port_b_first_bit_number = 5;
defparam ram_block1a69.port_b_last_address = 16383;
defparam ram_block1a69.port_b_logical_ram_depth = 16384;
defparam ram_block1a69.port_b_logical_ram_width = 64;
defparam ram_block1a69.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a69.port_b_read_enable_clock = "clock1";
defparam ram_block1a69.port_b_write_enable_clock = "clock1";
defparam ram_block1a69.ram_block_type = "auto";
defparam ram_block1a69.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a69.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a69.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a69.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a5(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[5]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.clk1_input_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "bidir_dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 13;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 8191;
defparam ram_block1a5.port_a_logical_ram_depth = 16384;
defparam ram_block1a5.port_a_logical_ram_width = 64;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 13;
defparam ram_block1a5.port_b_byte_enable_clock = "clock1";
defparam ram_block1a5.port_b_byte_enable_mask_width = 1;
defparam ram_block1a5.port_b_byte_size = 1;
defparam ram_block1a5.port_b_data_in_clock = "clock1";
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 8191;
defparam ram_block1a5.port_b_logical_ram_depth = 16384;
defparam ram_block1a5.port_b_logical_ram_width = 64;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.port_b_write_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a5.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a70(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[6]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a70_PORTADATAOUT_bus),
	.portbdataout(ram_block1a70_PORTBDATAOUT_bus));
defparam ram_block1a70.clk0_core_clock_enable = "ena0";
defparam ram_block1a70.clk0_input_clock_enable = "ena0";
defparam ram_block1a70.clk1_core_clock_enable = "ena1";
defparam ram_block1a70.clk1_input_clock_enable = "ena1";
defparam ram_block1a70.data_interleave_offset_in_bits = 1;
defparam ram_block1a70.data_interleave_width_in_bits = 1;
defparam ram_block1a70.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a70.init_file_layout = "port_a";
defparam ram_block1a70.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a70.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a70.operation_mode = "bidir_dual_port";
defparam ram_block1a70.port_a_address_clear = "none";
defparam ram_block1a70.port_a_address_width = 13;
defparam ram_block1a70.port_a_byte_enable_mask_width = 1;
defparam ram_block1a70.port_a_byte_size = 1;
defparam ram_block1a70.port_a_data_out_clear = "none";
defparam ram_block1a70.port_a_data_out_clock = "none";
defparam ram_block1a70.port_a_data_width = 1;
defparam ram_block1a70.port_a_first_address = 8192;
defparam ram_block1a70.port_a_first_bit_number = 6;
defparam ram_block1a70.port_a_last_address = 16383;
defparam ram_block1a70.port_a_logical_ram_depth = 16384;
defparam ram_block1a70.port_a_logical_ram_width = 64;
defparam ram_block1a70.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a70.port_b_address_clear = "none";
defparam ram_block1a70.port_b_address_clock = "clock1";
defparam ram_block1a70.port_b_address_width = 13;
defparam ram_block1a70.port_b_byte_enable_clock = "clock1";
defparam ram_block1a70.port_b_byte_enable_mask_width = 1;
defparam ram_block1a70.port_b_byte_size = 1;
defparam ram_block1a70.port_b_data_in_clock = "clock1";
defparam ram_block1a70.port_b_data_out_clear = "none";
defparam ram_block1a70.port_b_data_out_clock = "none";
defparam ram_block1a70.port_b_data_width = 1;
defparam ram_block1a70.port_b_first_address = 8192;
defparam ram_block1a70.port_b_first_bit_number = 6;
defparam ram_block1a70.port_b_last_address = 16383;
defparam ram_block1a70.port_b_logical_ram_depth = 16384;
defparam ram_block1a70.port_b_logical_ram_width = 64;
defparam ram_block1a70.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a70.port_b_read_enable_clock = "clock1";
defparam ram_block1a70.port_b_write_enable_clock = "clock1";
defparam ram_block1a70.ram_block_type = "auto";
defparam ram_block1a70.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a70.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a70.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a70.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a6(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[6]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.clk1_input_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "bidir_dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 13;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 8191;
defparam ram_block1a6.port_a_logical_ram_depth = 16384;
defparam ram_block1a6.port_a_logical_ram_width = 64;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 13;
defparam ram_block1a6.port_b_byte_enable_clock = "clock1";
defparam ram_block1a6.port_b_byte_enable_mask_width = 1;
defparam ram_block1a6.port_b_byte_size = 1;
defparam ram_block1a6.port_b_data_in_clock = "clock1";
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 8191;
defparam ram_block1a6.port_b_logical_ram_depth = 16384;
defparam ram_block1a6.port_b_logical_ram_width = 64;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.port_b_write_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a6.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a71(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[7]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a71_PORTADATAOUT_bus),
	.portbdataout(ram_block1a71_PORTBDATAOUT_bus));
defparam ram_block1a71.clk0_core_clock_enable = "ena0";
defparam ram_block1a71.clk0_input_clock_enable = "ena0";
defparam ram_block1a71.clk1_core_clock_enable = "ena1";
defparam ram_block1a71.clk1_input_clock_enable = "ena1";
defparam ram_block1a71.data_interleave_offset_in_bits = 1;
defparam ram_block1a71.data_interleave_width_in_bits = 1;
defparam ram_block1a71.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a71.init_file_layout = "port_a";
defparam ram_block1a71.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a71.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a71.operation_mode = "bidir_dual_port";
defparam ram_block1a71.port_a_address_clear = "none";
defparam ram_block1a71.port_a_address_width = 13;
defparam ram_block1a71.port_a_byte_enable_mask_width = 1;
defparam ram_block1a71.port_a_byte_size = 1;
defparam ram_block1a71.port_a_data_out_clear = "none";
defparam ram_block1a71.port_a_data_out_clock = "none";
defparam ram_block1a71.port_a_data_width = 1;
defparam ram_block1a71.port_a_first_address = 8192;
defparam ram_block1a71.port_a_first_bit_number = 7;
defparam ram_block1a71.port_a_last_address = 16383;
defparam ram_block1a71.port_a_logical_ram_depth = 16384;
defparam ram_block1a71.port_a_logical_ram_width = 64;
defparam ram_block1a71.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a71.port_b_address_clear = "none";
defparam ram_block1a71.port_b_address_clock = "clock1";
defparam ram_block1a71.port_b_address_width = 13;
defparam ram_block1a71.port_b_byte_enable_clock = "clock1";
defparam ram_block1a71.port_b_byte_enable_mask_width = 1;
defparam ram_block1a71.port_b_byte_size = 1;
defparam ram_block1a71.port_b_data_in_clock = "clock1";
defparam ram_block1a71.port_b_data_out_clear = "none";
defparam ram_block1a71.port_b_data_out_clock = "none";
defparam ram_block1a71.port_b_data_width = 1;
defparam ram_block1a71.port_b_first_address = 8192;
defparam ram_block1a71.port_b_first_bit_number = 7;
defparam ram_block1a71.port_b_last_address = 16383;
defparam ram_block1a71.port_b_logical_ram_depth = 16384;
defparam ram_block1a71.port_b_logical_ram_width = 64;
defparam ram_block1a71.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a71.port_b_read_enable_clock = "clock1";
defparam ram_block1a71.port_b_write_enable_clock = "clock1";
defparam ram_block1a71.ram_block_type = "auto";
defparam ram_block1a71.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a71.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a71.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a71.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a7(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[7]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[0]}),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.clk1_input_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "bidir_dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 13;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 8191;
defparam ram_block1a7.port_a_logical_ram_depth = 16384;
defparam ram_block1a7.port_a_logical_ram_width = 64;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 13;
defparam ram_block1a7.port_b_byte_enable_clock = "clock1";
defparam ram_block1a7.port_b_byte_enable_mask_width = 1;
defparam ram_block1a7.port_b_byte_size = 1;
defparam ram_block1a7.port_b_data_in_clock = "clock1";
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 8191;
defparam ram_block1a7.port_b_logical_ram_depth = 16384;
defparam ram_block1a7.port_b_logical_ram_width = 64;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.port_b_write_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a7.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a72(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[8]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a72_PORTADATAOUT_bus),
	.portbdataout(ram_block1a72_PORTBDATAOUT_bus));
defparam ram_block1a72.clk0_core_clock_enable = "ena0";
defparam ram_block1a72.clk0_input_clock_enable = "ena0";
defparam ram_block1a72.clk1_core_clock_enable = "ena1";
defparam ram_block1a72.clk1_input_clock_enable = "ena1";
defparam ram_block1a72.data_interleave_offset_in_bits = 1;
defparam ram_block1a72.data_interleave_width_in_bits = 1;
defparam ram_block1a72.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a72.init_file_layout = "port_a";
defparam ram_block1a72.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a72.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a72.operation_mode = "bidir_dual_port";
defparam ram_block1a72.port_a_address_clear = "none";
defparam ram_block1a72.port_a_address_width = 13;
defparam ram_block1a72.port_a_byte_enable_mask_width = 1;
defparam ram_block1a72.port_a_byte_size = 1;
defparam ram_block1a72.port_a_data_out_clear = "none";
defparam ram_block1a72.port_a_data_out_clock = "none";
defparam ram_block1a72.port_a_data_width = 1;
defparam ram_block1a72.port_a_first_address = 8192;
defparam ram_block1a72.port_a_first_bit_number = 8;
defparam ram_block1a72.port_a_last_address = 16383;
defparam ram_block1a72.port_a_logical_ram_depth = 16384;
defparam ram_block1a72.port_a_logical_ram_width = 64;
defparam ram_block1a72.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a72.port_b_address_clear = "none";
defparam ram_block1a72.port_b_address_clock = "clock1";
defparam ram_block1a72.port_b_address_width = 13;
defparam ram_block1a72.port_b_byte_enable_clock = "clock1";
defparam ram_block1a72.port_b_byte_enable_mask_width = 1;
defparam ram_block1a72.port_b_byte_size = 1;
defparam ram_block1a72.port_b_data_in_clock = "clock1";
defparam ram_block1a72.port_b_data_out_clear = "none";
defparam ram_block1a72.port_b_data_out_clock = "none";
defparam ram_block1a72.port_b_data_width = 1;
defparam ram_block1a72.port_b_first_address = 8192;
defparam ram_block1a72.port_b_first_bit_number = 8;
defparam ram_block1a72.port_b_last_address = 16383;
defparam ram_block1a72.port_b_logical_ram_depth = 16384;
defparam ram_block1a72.port_b_logical_ram_width = 64;
defparam ram_block1a72.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a72.port_b_read_enable_clock = "clock1";
defparam ram_block1a72.port_b_write_enable_clock = "clock1";
defparam ram_block1a72.ram_block_type = "auto";
defparam ram_block1a72.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a72.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a72.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a72.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a8(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[8]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.clk1_input_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "bidir_dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 13;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 8191;
defparam ram_block1a8.port_a_logical_ram_depth = 16384;
defparam ram_block1a8.port_a_logical_ram_width = 64;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 13;
defparam ram_block1a8.port_b_byte_enable_clock = "clock1";
defparam ram_block1a8.port_b_byte_enable_mask_width = 1;
defparam ram_block1a8.port_b_byte_size = 1;
defparam ram_block1a8.port_b_data_in_clock = "clock1";
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 8191;
defparam ram_block1a8.port_b_logical_ram_depth = 16384;
defparam ram_block1a8.port_b_logical_ram_width = 64;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.port_b_write_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a8.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a73(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[9]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a73_PORTADATAOUT_bus),
	.portbdataout(ram_block1a73_PORTBDATAOUT_bus));
defparam ram_block1a73.clk0_core_clock_enable = "ena0";
defparam ram_block1a73.clk0_input_clock_enable = "ena0";
defparam ram_block1a73.clk1_core_clock_enable = "ena1";
defparam ram_block1a73.clk1_input_clock_enable = "ena1";
defparam ram_block1a73.data_interleave_offset_in_bits = 1;
defparam ram_block1a73.data_interleave_width_in_bits = 1;
defparam ram_block1a73.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a73.init_file_layout = "port_a";
defparam ram_block1a73.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a73.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a73.operation_mode = "bidir_dual_port";
defparam ram_block1a73.port_a_address_clear = "none";
defparam ram_block1a73.port_a_address_width = 13;
defparam ram_block1a73.port_a_byte_enable_mask_width = 1;
defparam ram_block1a73.port_a_byte_size = 1;
defparam ram_block1a73.port_a_data_out_clear = "none";
defparam ram_block1a73.port_a_data_out_clock = "none";
defparam ram_block1a73.port_a_data_width = 1;
defparam ram_block1a73.port_a_first_address = 8192;
defparam ram_block1a73.port_a_first_bit_number = 9;
defparam ram_block1a73.port_a_last_address = 16383;
defparam ram_block1a73.port_a_logical_ram_depth = 16384;
defparam ram_block1a73.port_a_logical_ram_width = 64;
defparam ram_block1a73.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a73.port_b_address_clear = "none";
defparam ram_block1a73.port_b_address_clock = "clock1";
defparam ram_block1a73.port_b_address_width = 13;
defparam ram_block1a73.port_b_byte_enable_clock = "clock1";
defparam ram_block1a73.port_b_byte_enable_mask_width = 1;
defparam ram_block1a73.port_b_byte_size = 1;
defparam ram_block1a73.port_b_data_in_clock = "clock1";
defparam ram_block1a73.port_b_data_out_clear = "none";
defparam ram_block1a73.port_b_data_out_clock = "none";
defparam ram_block1a73.port_b_data_width = 1;
defparam ram_block1a73.port_b_first_address = 8192;
defparam ram_block1a73.port_b_first_bit_number = 9;
defparam ram_block1a73.port_b_last_address = 16383;
defparam ram_block1a73.port_b_logical_ram_depth = 16384;
defparam ram_block1a73.port_b_logical_ram_width = 64;
defparam ram_block1a73.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a73.port_b_read_enable_clock = "clock1";
defparam ram_block1a73.port_b_write_enable_clock = "clock1";
defparam ram_block1a73.ram_block_type = "auto";
defparam ram_block1a73.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a73.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a73.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a73.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a9(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[9]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.clk1_input_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "bidir_dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 13;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 8191;
defparam ram_block1a9.port_a_logical_ram_depth = 16384;
defparam ram_block1a9.port_a_logical_ram_width = 64;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 13;
defparam ram_block1a9.port_b_byte_enable_clock = "clock1";
defparam ram_block1a9.port_b_byte_enable_mask_width = 1;
defparam ram_block1a9.port_b_byte_size = 1;
defparam ram_block1a9.port_b_data_in_clock = "clock1";
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 8191;
defparam ram_block1a9.port_b_logical_ram_depth = 16384;
defparam ram_block1a9.port_b_logical_ram_width = 64;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.port_b_write_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a9.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a74(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[10]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a74_PORTADATAOUT_bus),
	.portbdataout(ram_block1a74_PORTBDATAOUT_bus));
defparam ram_block1a74.clk0_core_clock_enable = "ena0";
defparam ram_block1a74.clk0_input_clock_enable = "ena0";
defparam ram_block1a74.clk1_core_clock_enable = "ena1";
defparam ram_block1a74.clk1_input_clock_enable = "ena1";
defparam ram_block1a74.data_interleave_offset_in_bits = 1;
defparam ram_block1a74.data_interleave_width_in_bits = 1;
defparam ram_block1a74.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a74.init_file_layout = "port_a";
defparam ram_block1a74.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a74.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a74.operation_mode = "bidir_dual_port";
defparam ram_block1a74.port_a_address_clear = "none";
defparam ram_block1a74.port_a_address_width = 13;
defparam ram_block1a74.port_a_byte_enable_mask_width = 1;
defparam ram_block1a74.port_a_byte_size = 1;
defparam ram_block1a74.port_a_data_out_clear = "none";
defparam ram_block1a74.port_a_data_out_clock = "none";
defparam ram_block1a74.port_a_data_width = 1;
defparam ram_block1a74.port_a_first_address = 8192;
defparam ram_block1a74.port_a_first_bit_number = 10;
defparam ram_block1a74.port_a_last_address = 16383;
defparam ram_block1a74.port_a_logical_ram_depth = 16384;
defparam ram_block1a74.port_a_logical_ram_width = 64;
defparam ram_block1a74.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a74.port_b_address_clear = "none";
defparam ram_block1a74.port_b_address_clock = "clock1";
defparam ram_block1a74.port_b_address_width = 13;
defparam ram_block1a74.port_b_byte_enable_clock = "clock1";
defparam ram_block1a74.port_b_byte_enable_mask_width = 1;
defparam ram_block1a74.port_b_byte_size = 1;
defparam ram_block1a74.port_b_data_in_clock = "clock1";
defparam ram_block1a74.port_b_data_out_clear = "none";
defparam ram_block1a74.port_b_data_out_clock = "none";
defparam ram_block1a74.port_b_data_width = 1;
defparam ram_block1a74.port_b_first_address = 8192;
defparam ram_block1a74.port_b_first_bit_number = 10;
defparam ram_block1a74.port_b_last_address = 16383;
defparam ram_block1a74.port_b_logical_ram_depth = 16384;
defparam ram_block1a74.port_b_logical_ram_width = 64;
defparam ram_block1a74.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a74.port_b_read_enable_clock = "clock1";
defparam ram_block1a74.port_b_write_enable_clock = "clock1";
defparam ram_block1a74.ram_block_type = "auto";
defparam ram_block1a74.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a74.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a74.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a74.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a10(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[10]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.clk1_input_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "bidir_dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 13;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 8191;
defparam ram_block1a10.port_a_logical_ram_depth = 16384;
defparam ram_block1a10.port_a_logical_ram_width = 64;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 13;
defparam ram_block1a10.port_b_byte_enable_clock = "clock1";
defparam ram_block1a10.port_b_byte_enable_mask_width = 1;
defparam ram_block1a10.port_b_byte_size = 1;
defparam ram_block1a10.port_b_data_in_clock = "clock1";
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 8191;
defparam ram_block1a10.port_b_logical_ram_depth = 16384;
defparam ram_block1a10.port_b_logical_ram_width = 64;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.port_b_write_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a10.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a75(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[11]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a75_PORTADATAOUT_bus),
	.portbdataout(ram_block1a75_PORTBDATAOUT_bus));
defparam ram_block1a75.clk0_core_clock_enable = "ena0";
defparam ram_block1a75.clk0_input_clock_enable = "ena0";
defparam ram_block1a75.clk1_core_clock_enable = "ena1";
defparam ram_block1a75.clk1_input_clock_enable = "ena1";
defparam ram_block1a75.data_interleave_offset_in_bits = 1;
defparam ram_block1a75.data_interleave_width_in_bits = 1;
defparam ram_block1a75.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a75.init_file_layout = "port_a";
defparam ram_block1a75.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a75.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a75.operation_mode = "bidir_dual_port";
defparam ram_block1a75.port_a_address_clear = "none";
defparam ram_block1a75.port_a_address_width = 13;
defparam ram_block1a75.port_a_byte_enable_mask_width = 1;
defparam ram_block1a75.port_a_byte_size = 1;
defparam ram_block1a75.port_a_data_out_clear = "none";
defparam ram_block1a75.port_a_data_out_clock = "none";
defparam ram_block1a75.port_a_data_width = 1;
defparam ram_block1a75.port_a_first_address = 8192;
defparam ram_block1a75.port_a_first_bit_number = 11;
defparam ram_block1a75.port_a_last_address = 16383;
defparam ram_block1a75.port_a_logical_ram_depth = 16384;
defparam ram_block1a75.port_a_logical_ram_width = 64;
defparam ram_block1a75.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a75.port_b_address_clear = "none";
defparam ram_block1a75.port_b_address_clock = "clock1";
defparam ram_block1a75.port_b_address_width = 13;
defparam ram_block1a75.port_b_byte_enable_clock = "clock1";
defparam ram_block1a75.port_b_byte_enable_mask_width = 1;
defparam ram_block1a75.port_b_byte_size = 1;
defparam ram_block1a75.port_b_data_in_clock = "clock1";
defparam ram_block1a75.port_b_data_out_clear = "none";
defparam ram_block1a75.port_b_data_out_clock = "none";
defparam ram_block1a75.port_b_data_width = 1;
defparam ram_block1a75.port_b_first_address = 8192;
defparam ram_block1a75.port_b_first_bit_number = 11;
defparam ram_block1a75.port_b_last_address = 16383;
defparam ram_block1a75.port_b_logical_ram_depth = 16384;
defparam ram_block1a75.port_b_logical_ram_width = 64;
defparam ram_block1a75.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a75.port_b_read_enable_clock = "clock1";
defparam ram_block1a75.port_b_write_enable_clock = "clock1";
defparam ram_block1a75.ram_block_type = "auto";
defparam ram_block1a75.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a75.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a75.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a75.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a11(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[11]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.clk1_input_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "bidir_dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 13;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 8191;
defparam ram_block1a11.port_a_logical_ram_depth = 16384;
defparam ram_block1a11.port_a_logical_ram_width = 64;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 13;
defparam ram_block1a11.port_b_byte_enable_clock = "clock1";
defparam ram_block1a11.port_b_byte_enable_mask_width = 1;
defparam ram_block1a11.port_b_byte_size = 1;
defparam ram_block1a11.port_b_data_in_clock = "clock1";
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 8191;
defparam ram_block1a11.port_b_logical_ram_depth = 16384;
defparam ram_block1a11.port_b_logical_ram_width = 64;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.port_b_write_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a11.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a76(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[12]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a76_PORTADATAOUT_bus),
	.portbdataout(ram_block1a76_PORTBDATAOUT_bus));
defparam ram_block1a76.clk0_core_clock_enable = "ena0";
defparam ram_block1a76.clk0_input_clock_enable = "ena0";
defparam ram_block1a76.clk1_core_clock_enable = "ena1";
defparam ram_block1a76.clk1_input_clock_enable = "ena1";
defparam ram_block1a76.data_interleave_offset_in_bits = 1;
defparam ram_block1a76.data_interleave_width_in_bits = 1;
defparam ram_block1a76.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a76.init_file_layout = "port_a";
defparam ram_block1a76.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a76.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a76.operation_mode = "bidir_dual_port";
defparam ram_block1a76.port_a_address_clear = "none";
defparam ram_block1a76.port_a_address_width = 13;
defparam ram_block1a76.port_a_byte_enable_mask_width = 1;
defparam ram_block1a76.port_a_byte_size = 1;
defparam ram_block1a76.port_a_data_out_clear = "none";
defparam ram_block1a76.port_a_data_out_clock = "none";
defparam ram_block1a76.port_a_data_width = 1;
defparam ram_block1a76.port_a_first_address = 8192;
defparam ram_block1a76.port_a_first_bit_number = 12;
defparam ram_block1a76.port_a_last_address = 16383;
defparam ram_block1a76.port_a_logical_ram_depth = 16384;
defparam ram_block1a76.port_a_logical_ram_width = 64;
defparam ram_block1a76.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a76.port_b_address_clear = "none";
defparam ram_block1a76.port_b_address_clock = "clock1";
defparam ram_block1a76.port_b_address_width = 13;
defparam ram_block1a76.port_b_byte_enable_clock = "clock1";
defparam ram_block1a76.port_b_byte_enable_mask_width = 1;
defparam ram_block1a76.port_b_byte_size = 1;
defparam ram_block1a76.port_b_data_in_clock = "clock1";
defparam ram_block1a76.port_b_data_out_clear = "none";
defparam ram_block1a76.port_b_data_out_clock = "none";
defparam ram_block1a76.port_b_data_width = 1;
defparam ram_block1a76.port_b_first_address = 8192;
defparam ram_block1a76.port_b_first_bit_number = 12;
defparam ram_block1a76.port_b_last_address = 16383;
defparam ram_block1a76.port_b_logical_ram_depth = 16384;
defparam ram_block1a76.port_b_logical_ram_width = 64;
defparam ram_block1a76.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a76.port_b_read_enable_clock = "clock1";
defparam ram_block1a76.port_b_write_enable_clock = "clock1";
defparam ram_block1a76.ram_block_type = "auto";
defparam ram_block1a76.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a76.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a76.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a76.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a12(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[12]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.clk1_input_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "bidir_dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 13;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 8191;
defparam ram_block1a12.port_a_logical_ram_depth = 16384;
defparam ram_block1a12.port_a_logical_ram_width = 64;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 13;
defparam ram_block1a12.port_b_byte_enable_clock = "clock1";
defparam ram_block1a12.port_b_byte_enable_mask_width = 1;
defparam ram_block1a12.port_b_byte_size = 1;
defparam ram_block1a12.port_b_data_in_clock = "clock1";
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 8191;
defparam ram_block1a12.port_b_logical_ram_depth = 16384;
defparam ram_block1a12.port_b_logical_ram_width = 64;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.port_b_write_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a12.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a77(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[13]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a77_PORTADATAOUT_bus),
	.portbdataout(ram_block1a77_PORTBDATAOUT_bus));
defparam ram_block1a77.clk0_core_clock_enable = "ena0";
defparam ram_block1a77.clk0_input_clock_enable = "ena0";
defparam ram_block1a77.clk1_core_clock_enable = "ena1";
defparam ram_block1a77.clk1_input_clock_enable = "ena1";
defparam ram_block1a77.data_interleave_offset_in_bits = 1;
defparam ram_block1a77.data_interleave_width_in_bits = 1;
defparam ram_block1a77.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a77.init_file_layout = "port_a";
defparam ram_block1a77.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a77.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a77.operation_mode = "bidir_dual_port";
defparam ram_block1a77.port_a_address_clear = "none";
defparam ram_block1a77.port_a_address_width = 13;
defparam ram_block1a77.port_a_byte_enable_mask_width = 1;
defparam ram_block1a77.port_a_byte_size = 1;
defparam ram_block1a77.port_a_data_out_clear = "none";
defparam ram_block1a77.port_a_data_out_clock = "none";
defparam ram_block1a77.port_a_data_width = 1;
defparam ram_block1a77.port_a_first_address = 8192;
defparam ram_block1a77.port_a_first_bit_number = 13;
defparam ram_block1a77.port_a_last_address = 16383;
defparam ram_block1a77.port_a_logical_ram_depth = 16384;
defparam ram_block1a77.port_a_logical_ram_width = 64;
defparam ram_block1a77.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a77.port_b_address_clear = "none";
defparam ram_block1a77.port_b_address_clock = "clock1";
defparam ram_block1a77.port_b_address_width = 13;
defparam ram_block1a77.port_b_byte_enable_clock = "clock1";
defparam ram_block1a77.port_b_byte_enable_mask_width = 1;
defparam ram_block1a77.port_b_byte_size = 1;
defparam ram_block1a77.port_b_data_in_clock = "clock1";
defparam ram_block1a77.port_b_data_out_clear = "none";
defparam ram_block1a77.port_b_data_out_clock = "none";
defparam ram_block1a77.port_b_data_width = 1;
defparam ram_block1a77.port_b_first_address = 8192;
defparam ram_block1a77.port_b_first_bit_number = 13;
defparam ram_block1a77.port_b_last_address = 16383;
defparam ram_block1a77.port_b_logical_ram_depth = 16384;
defparam ram_block1a77.port_b_logical_ram_width = 64;
defparam ram_block1a77.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a77.port_b_read_enable_clock = "clock1";
defparam ram_block1a77.port_b_write_enable_clock = "clock1";
defparam ram_block1a77.ram_block_type = "auto";
defparam ram_block1a77.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a77.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a77.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a77.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a13(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[13]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.clk1_input_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "bidir_dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 13;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 8191;
defparam ram_block1a13.port_a_logical_ram_depth = 16384;
defparam ram_block1a13.port_a_logical_ram_width = 64;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 13;
defparam ram_block1a13.port_b_byte_enable_clock = "clock1";
defparam ram_block1a13.port_b_byte_enable_mask_width = 1;
defparam ram_block1a13.port_b_byte_size = 1;
defparam ram_block1a13.port_b_data_in_clock = "clock1";
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 8191;
defparam ram_block1a13.port_b_logical_ram_depth = 16384;
defparam ram_block1a13.port_b_logical_ram_width = 64;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.port_b_write_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a13.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a78(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[14]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a78_PORTADATAOUT_bus),
	.portbdataout(ram_block1a78_PORTBDATAOUT_bus));
defparam ram_block1a78.clk0_core_clock_enable = "ena0";
defparam ram_block1a78.clk0_input_clock_enable = "ena0";
defparam ram_block1a78.clk1_core_clock_enable = "ena1";
defparam ram_block1a78.clk1_input_clock_enable = "ena1";
defparam ram_block1a78.data_interleave_offset_in_bits = 1;
defparam ram_block1a78.data_interleave_width_in_bits = 1;
defparam ram_block1a78.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a78.init_file_layout = "port_a";
defparam ram_block1a78.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a78.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a78.operation_mode = "bidir_dual_port";
defparam ram_block1a78.port_a_address_clear = "none";
defparam ram_block1a78.port_a_address_width = 13;
defparam ram_block1a78.port_a_byte_enable_mask_width = 1;
defparam ram_block1a78.port_a_byte_size = 1;
defparam ram_block1a78.port_a_data_out_clear = "none";
defparam ram_block1a78.port_a_data_out_clock = "none";
defparam ram_block1a78.port_a_data_width = 1;
defparam ram_block1a78.port_a_first_address = 8192;
defparam ram_block1a78.port_a_first_bit_number = 14;
defparam ram_block1a78.port_a_last_address = 16383;
defparam ram_block1a78.port_a_logical_ram_depth = 16384;
defparam ram_block1a78.port_a_logical_ram_width = 64;
defparam ram_block1a78.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a78.port_b_address_clear = "none";
defparam ram_block1a78.port_b_address_clock = "clock1";
defparam ram_block1a78.port_b_address_width = 13;
defparam ram_block1a78.port_b_byte_enable_clock = "clock1";
defparam ram_block1a78.port_b_byte_enable_mask_width = 1;
defparam ram_block1a78.port_b_byte_size = 1;
defparam ram_block1a78.port_b_data_in_clock = "clock1";
defparam ram_block1a78.port_b_data_out_clear = "none";
defparam ram_block1a78.port_b_data_out_clock = "none";
defparam ram_block1a78.port_b_data_width = 1;
defparam ram_block1a78.port_b_first_address = 8192;
defparam ram_block1a78.port_b_first_bit_number = 14;
defparam ram_block1a78.port_b_last_address = 16383;
defparam ram_block1a78.port_b_logical_ram_depth = 16384;
defparam ram_block1a78.port_b_logical_ram_width = 64;
defparam ram_block1a78.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a78.port_b_read_enable_clock = "clock1";
defparam ram_block1a78.port_b_write_enable_clock = "clock1";
defparam ram_block1a78.ram_block_type = "auto";
defparam ram_block1a78.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a78.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a78.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a78.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a14(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[14]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.clk1_input_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "bidir_dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 13;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 8191;
defparam ram_block1a14.port_a_logical_ram_depth = 16384;
defparam ram_block1a14.port_a_logical_ram_width = 64;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 13;
defparam ram_block1a14.port_b_byte_enable_clock = "clock1";
defparam ram_block1a14.port_b_byte_enable_mask_width = 1;
defparam ram_block1a14.port_b_byte_size = 1;
defparam ram_block1a14.port_b_data_in_clock = "clock1";
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 8191;
defparam ram_block1a14.port_b_logical_ram_depth = 16384;
defparam ram_block1a14.port_b_logical_ram_width = 64;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.port_b_write_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a14.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a79(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[15]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a79_PORTADATAOUT_bus),
	.portbdataout(ram_block1a79_PORTBDATAOUT_bus));
defparam ram_block1a79.clk0_core_clock_enable = "ena0";
defparam ram_block1a79.clk0_input_clock_enable = "ena0";
defparam ram_block1a79.clk1_core_clock_enable = "ena1";
defparam ram_block1a79.clk1_input_clock_enable = "ena1";
defparam ram_block1a79.data_interleave_offset_in_bits = 1;
defparam ram_block1a79.data_interleave_width_in_bits = 1;
defparam ram_block1a79.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a79.init_file_layout = "port_a";
defparam ram_block1a79.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a79.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a79.operation_mode = "bidir_dual_port";
defparam ram_block1a79.port_a_address_clear = "none";
defparam ram_block1a79.port_a_address_width = 13;
defparam ram_block1a79.port_a_byte_enable_mask_width = 1;
defparam ram_block1a79.port_a_byte_size = 1;
defparam ram_block1a79.port_a_data_out_clear = "none";
defparam ram_block1a79.port_a_data_out_clock = "none";
defparam ram_block1a79.port_a_data_width = 1;
defparam ram_block1a79.port_a_first_address = 8192;
defparam ram_block1a79.port_a_first_bit_number = 15;
defparam ram_block1a79.port_a_last_address = 16383;
defparam ram_block1a79.port_a_logical_ram_depth = 16384;
defparam ram_block1a79.port_a_logical_ram_width = 64;
defparam ram_block1a79.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a79.port_b_address_clear = "none";
defparam ram_block1a79.port_b_address_clock = "clock1";
defparam ram_block1a79.port_b_address_width = 13;
defparam ram_block1a79.port_b_byte_enable_clock = "clock1";
defparam ram_block1a79.port_b_byte_enable_mask_width = 1;
defparam ram_block1a79.port_b_byte_size = 1;
defparam ram_block1a79.port_b_data_in_clock = "clock1";
defparam ram_block1a79.port_b_data_out_clear = "none";
defparam ram_block1a79.port_b_data_out_clock = "none";
defparam ram_block1a79.port_b_data_width = 1;
defparam ram_block1a79.port_b_first_address = 8192;
defparam ram_block1a79.port_b_first_bit_number = 15;
defparam ram_block1a79.port_b_last_address = 16383;
defparam ram_block1a79.port_b_logical_ram_depth = 16384;
defparam ram_block1a79.port_b_logical_ram_width = 64;
defparam ram_block1a79.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a79.port_b_read_enable_clock = "clock1";
defparam ram_block1a79.port_b_write_enable_clock = "clock1";
defparam ram_block1a79.ram_block_type = "auto";
defparam ram_block1a79.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a79.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a79.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a79.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a15(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[15]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[1]}),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.clk1_input_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "bidir_dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 13;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 8191;
defparam ram_block1a15.port_a_logical_ram_depth = 16384;
defparam ram_block1a15.port_a_logical_ram_width = 64;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 13;
defparam ram_block1a15.port_b_byte_enable_clock = "clock1";
defparam ram_block1a15.port_b_byte_enable_mask_width = 1;
defparam ram_block1a15.port_b_byte_size = 1;
defparam ram_block1a15.port_b_data_in_clock = "clock1";
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 8191;
defparam ram_block1a15.port_b_logical_ram_depth = 16384;
defparam ram_block1a15.port_b_logical_ram_width = 64;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.port_b_write_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a15.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a80(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[16]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a80_PORTADATAOUT_bus),
	.portbdataout(ram_block1a80_PORTBDATAOUT_bus));
defparam ram_block1a80.clk0_core_clock_enable = "ena0";
defparam ram_block1a80.clk0_input_clock_enable = "ena0";
defparam ram_block1a80.clk1_core_clock_enable = "ena1";
defparam ram_block1a80.clk1_input_clock_enable = "ena1";
defparam ram_block1a80.data_interleave_offset_in_bits = 1;
defparam ram_block1a80.data_interleave_width_in_bits = 1;
defparam ram_block1a80.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a80.init_file_layout = "port_a";
defparam ram_block1a80.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a80.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a80.operation_mode = "bidir_dual_port";
defparam ram_block1a80.port_a_address_clear = "none";
defparam ram_block1a80.port_a_address_width = 13;
defparam ram_block1a80.port_a_byte_enable_mask_width = 1;
defparam ram_block1a80.port_a_byte_size = 1;
defparam ram_block1a80.port_a_data_out_clear = "none";
defparam ram_block1a80.port_a_data_out_clock = "none";
defparam ram_block1a80.port_a_data_width = 1;
defparam ram_block1a80.port_a_first_address = 8192;
defparam ram_block1a80.port_a_first_bit_number = 16;
defparam ram_block1a80.port_a_last_address = 16383;
defparam ram_block1a80.port_a_logical_ram_depth = 16384;
defparam ram_block1a80.port_a_logical_ram_width = 64;
defparam ram_block1a80.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a80.port_b_address_clear = "none";
defparam ram_block1a80.port_b_address_clock = "clock1";
defparam ram_block1a80.port_b_address_width = 13;
defparam ram_block1a80.port_b_byte_enable_clock = "clock1";
defparam ram_block1a80.port_b_byte_enable_mask_width = 1;
defparam ram_block1a80.port_b_byte_size = 1;
defparam ram_block1a80.port_b_data_in_clock = "clock1";
defparam ram_block1a80.port_b_data_out_clear = "none";
defparam ram_block1a80.port_b_data_out_clock = "none";
defparam ram_block1a80.port_b_data_width = 1;
defparam ram_block1a80.port_b_first_address = 8192;
defparam ram_block1a80.port_b_first_bit_number = 16;
defparam ram_block1a80.port_b_last_address = 16383;
defparam ram_block1a80.port_b_logical_ram_depth = 16384;
defparam ram_block1a80.port_b_logical_ram_width = 64;
defparam ram_block1a80.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a80.port_b_read_enable_clock = "clock1";
defparam ram_block1a80.port_b_write_enable_clock = "clock1";
defparam ram_block1a80.ram_block_type = "auto";
defparam ram_block1a80.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a80.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a80.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a80.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a16(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[16]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus));
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.clk1_core_clock_enable = "ena1";
defparam ram_block1a16.clk1_input_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "bidir_dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 13;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 8191;
defparam ram_block1a16.port_a_logical_ram_depth = 16384;
defparam ram_block1a16.port_a_logical_ram_width = 64;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 13;
defparam ram_block1a16.port_b_byte_enable_clock = "clock1";
defparam ram_block1a16.port_b_byte_enable_mask_width = 1;
defparam ram_block1a16.port_b_byte_size = 1;
defparam ram_block1a16.port_b_data_in_clock = "clock1";
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 8191;
defparam ram_block1a16.port_b_logical_ram_depth = 16384;
defparam ram_block1a16.port_b_logical_ram_width = 64;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.port_b_write_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a16.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a81(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[17]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a81_PORTADATAOUT_bus),
	.portbdataout(ram_block1a81_PORTBDATAOUT_bus));
defparam ram_block1a81.clk0_core_clock_enable = "ena0";
defparam ram_block1a81.clk0_input_clock_enable = "ena0";
defparam ram_block1a81.clk1_core_clock_enable = "ena1";
defparam ram_block1a81.clk1_input_clock_enable = "ena1";
defparam ram_block1a81.data_interleave_offset_in_bits = 1;
defparam ram_block1a81.data_interleave_width_in_bits = 1;
defparam ram_block1a81.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a81.init_file_layout = "port_a";
defparam ram_block1a81.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a81.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a81.operation_mode = "bidir_dual_port";
defparam ram_block1a81.port_a_address_clear = "none";
defparam ram_block1a81.port_a_address_width = 13;
defparam ram_block1a81.port_a_byte_enable_mask_width = 1;
defparam ram_block1a81.port_a_byte_size = 1;
defparam ram_block1a81.port_a_data_out_clear = "none";
defparam ram_block1a81.port_a_data_out_clock = "none";
defparam ram_block1a81.port_a_data_width = 1;
defparam ram_block1a81.port_a_first_address = 8192;
defparam ram_block1a81.port_a_first_bit_number = 17;
defparam ram_block1a81.port_a_last_address = 16383;
defparam ram_block1a81.port_a_logical_ram_depth = 16384;
defparam ram_block1a81.port_a_logical_ram_width = 64;
defparam ram_block1a81.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a81.port_b_address_clear = "none";
defparam ram_block1a81.port_b_address_clock = "clock1";
defparam ram_block1a81.port_b_address_width = 13;
defparam ram_block1a81.port_b_byte_enable_clock = "clock1";
defparam ram_block1a81.port_b_byte_enable_mask_width = 1;
defparam ram_block1a81.port_b_byte_size = 1;
defparam ram_block1a81.port_b_data_in_clock = "clock1";
defparam ram_block1a81.port_b_data_out_clear = "none";
defparam ram_block1a81.port_b_data_out_clock = "none";
defparam ram_block1a81.port_b_data_width = 1;
defparam ram_block1a81.port_b_first_address = 8192;
defparam ram_block1a81.port_b_first_bit_number = 17;
defparam ram_block1a81.port_b_last_address = 16383;
defparam ram_block1a81.port_b_logical_ram_depth = 16384;
defparam ram_block1a81.port_b_logical_ram_width = 64;
defparam ram_block1a81.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a81.port_b_read_enable_clock = "clock1";
defparam ram_block1a81.port_b_write_enable_clock = "clock1";
defparam ram_block1a81.ram_block_type = "auto";
defparam ram_block1a81.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a81.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a81.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a81.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a17(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[17]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus));
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.clk1_core_clock_enable = "ena1";
defparam ram_block1a17.clk1_input_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "bidir_dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 13;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 8191;
defparam ram_block1a17.port_a_logical_ram_depth = 16384;
defparam ram_block1a17.port_a_logical_ram_width = 64;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 13;
defparam ram_block1a17.port_b_byte_enable_clock = "clock1";
defparam ram_block1a17.port_b_byte_enable_mask_width = 1;
defparam ram_block1a17.port_b_byte_size = 1;
defparam ram_block1a17.port_b_data_in_clock = "clock1";
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 8191;
defparam ram_block1a17.port_b_logical_ram_depth = 16384;
defparam ram_block1a17.port_b_logical_ram_width = 64;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.port_b_write_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a17.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a82(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[18]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a82_PORTADATAOUT_bus),
	.portbdataout(ram_block1a82_PORTBDATAOUT_bus));
defparam ram_block1a82.clk0_core_clock_enable = "ena0";
defparam ram_block1a82.clk0_input_clock_enable = "ena0";
defparam ram_block1a82.clk1_core_clock_enable = "ena1";
defparam ram_block1a82.clk1_input_clock_enable = "ena1";
defparam ram_block1a82.data_interleave_offset_in_bits = 1;
defparam ram_block1a82.data_interleave_width_in_bits = 1;
defparam ram_block1a82.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a82.init_file_layout = "port_a";
defparam ram_block1a82.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a82.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a82.operation_mode = "bidir_dual_port";
defparam ram_block1a82.port_a_address_clear = "none";
defparam ram_block1a82.port_a_address_width = 13;
defparam ram_block1a82.port_a_byte_enable_mask_width = 1;
defparam ram_block1a82.port_a_byte_size = 1;
defparam ram_block1a82.port_a_data_out_clear = "none";
defparam ram_block1a82.port_a_data_out_clock = "none";
defparam ram_block1a82.port_a_data_width = 1;
defparam ram_block1a82.port_a_first_address = 8192;
defparam ram_block1a82.port_a_first_bit_number = 18;
defparam ram_block1a82.port_a_last_address = 16383;
defparam ram_block1a82.port_a_logical_ram_depth = 16384;
defparam ram_block1a82.port_a_logical_ram_width = 64;
defparam ram_block1a82.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a82.port_b_address_clear = "none";
defparam ram_block1a82.port_b_address_clock = "clock1";
defparam ram_block1a82.port_b_address_width = 13;
defparam ram_block1a82.port_b_byte_enable_clock = "clock1";
defparam ram_block1a82.port_b_byte_enable_mask_width = 1;
defparam ram_block1a82.port_b_byte_size = 1;
defparam ram_block1a82.port_b_data_in_clock = "clock1";
defparam ram_block1a82.port_b_data_out_clear = "none";
defparam ram_block1a82.port_b_data_out_clock = "none";
defparam ram_block1a82.port_b_data_width = 1;
defparam ram_block1a82.port_b_first_address = 8192;
defparam ram_block1a82.port_b_first_bit_number = 18;
defparam ram_block1a82.port_b_last_address = 16383;
defparam ram_block1a82.port_b_logical_ram_depth = 16384;
defparam ram_block1a82.port_b_logical_ram_width = 64;
defparam ram_block1a82.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a82.port_b_read_enable_clock = "clock1";
defparam ram_block1a82.port_b_write_enable_clock = "clock1";
defparam ram_block1a82.ram_block_type = "auto";
defparam ram_block1a82.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a82.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a82.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a82.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a18(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[18]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus));
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.clk1_core_clock_enable = "ena1";
defparam ram_block1a18.clk1_input_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "bidir_dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 13;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 8191;
defparam ram_block1a18.port_a_logical_ram_depth = 16384;
defparam ram_block1a18.port_a_logical_ram_width = 64;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 13;
defparam ram_block1a18.port_b_byte_enable_clock = "clock1";
defparam ram_block1a18.port_b_byte_enable_mask_width = 1;
defparam ram_block1a18.port_b_byte_size = 1;
defparam ram_block1a18.port_b_data_in_clock = "clock1";
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 8191;
defparam ram_block1a18.port_b_logical_ram_depth = 16384;
defparam ram_block1a18.port_b_logical_ram_width = 64;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.port_b_write_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a18.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a83(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[19]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a83_PORTADATAOUT_bus),
	.portbdataout(ram_block1a83_PORTBDATAOUT_bus));
defparam ram_block1a83.clk0_core_clock_enable = "ena0";
defparam ram_block1a83.clk0_input_clock_enable = "ena0";
defparam ram_block1a83.clk1_core_clock_enable = "ena1";
defparam ram_block1a83.clk1_input_clock_enable = "ena1";
defparam ram_block1a83.data_interleave_offset_in_bits = 1;
defparam ram_block1a83.data_interleave_width_in_bits = 1;
defparam ram_block1a83.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a83.init_file_layout = "port_a";
defparam ram_block1a83.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a83.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a83.operation_mode = "bidir_dual_port";
defparam ram_block1a83.port_a_address_clear = "none";
defparam ram_block1a83.port_a_address_width = 13;
defparam ram_block1a83.port_a_byte_enable_mask_width = 1;
defparam ram_block1a83.port_a_byte_size = 1;
defparam ram_block1a83.port_a_data_out_clear = "none";
defparam ram_block1a83.port_a_data_out_clock = "none";
defparam ram_block1a83.port_a_data_width = 1;
defparam ram_block1a83.port_a_first_address = 8192;
defparam ram_block1a83.port_a_first_bit_number = 19;
defparam ram_block1a83.port_a_last_address = 16383;
defparam ram_block1a83.port_a_logical_ram_depth = 16384;
defparam ram_block1a83.port_a_logical_ram_width = 64;
defparam ram_block1a83.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a83.port_b_address_clear = "none";
defparam ram_block1a83.port_b_address_clock = "clock1";
defparam ram_block1a83.port_b_address_width = 13;
defparam ram_block1a83.port_b_byte_enable_clock = "clock1";
defparam ram_block1a83.port_b_byte_enable_mask_width = 1;
defparam ram_block1a83.port_b_byte_size = 1;
defparam ram_block1a83.port_b_data_in_clock = "clock1";
defparam ram_block1a83.port_b_data_out_clear = "none";
defparam ram_block1a83.port_b_data_out_clock = "none";
defparam ram_block1a83.port_b_data_width = 1;
defparam ram_block1a83.port_b_first_address = 8192;
defparam ram_block1a83.port_b_first_bit_number = 19;
defparam ram_block1a83.port_b_last_address = 16383;
defparam ram_block1a83.port_b_logical_ram_depth = 16384;
defparam ram_block1a83.port_b_logical_ram_width = 64;
defparam ram_block1a83.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a83.port_b_read_enable_clock = "clock1";
defparam ram_block1a83.port_b_write_enable_clock = "clock1";
defparam ram_block1a83.ram_block_type = "auto";
defparam ram_block1a83.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a83.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a83.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a83.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a19(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[19]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus));
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.clk1_core_clock_enable = "ena1";
defparam ram_block1a19.clk1_input_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "bidir_dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 13;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 8191;
defparam ram_block1a19.port_a_logical_ram_depth = 16384;
defparam ram_block1a19.port_a_logical_ram_width = 64;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 13;
defparam ram_block1a19.port_b_byte_enable_clock = "clock1";
defparam ram_block1a19.port_b_byte_enable_mask_width = 1;
defparam ram_block1a19.port_b_byte_size = 1;
defparam ram_block1a19.port_b_data_in_clock = "clock1";
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 8191;
defparam ram_block1a19.port_b_logical_ram_depth = 16384;
defparam ram_block1a19.port_b_logical_ram_width = 64;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.port_b_write_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a19.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a84(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[20]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a84_PORTADATAOUT_bus),
	.portbdataout(ram_block1a84_PORTBDATAOUT_bus));
defparam ram_block1a84.clk0_core_clock_enable = "ena0";
defparam ram_block1a84.clk0_input_clock_enable = "ena0";
defparam ram_block1a84.clk1_core_clock_enable = "ena1";
defparam ram_block1a84.clk1_input_clock_enable = "ena1";
defparam ram_block1a84.data_interleave_offset_in_bits = 1;
defparam ram_block1a84.data_interleave_width_in_bits = 1;
defparam ram_block1a84.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a84.init_file_layout = "port_a";
defparam ram_block1a84.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a84.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a84.operation_mode = "bidir_dual_port";
defparam ram_block1a84.port_a_address_clear = "none";
defparam ram_block1a84.port_a_address_width = 13;
defparam ram_block1a84.port_a_byte_enable_mask_width = 1;
defparam ram_block1a84.port_a_byte_size = 1;
defparam ram_block1a84.port_a_data_out_clear = "none";
defparam ram_block1a84.port_a_data_out_clock = "none";
defparam ram_block1a84.port_a_data_width = 1;
defparam ram_block1a84.port_a_first_address = 8192;
defparam ram_block1a84.port_a_first_bit_number = 20;
defparam ram_block1a84.port_a_last_address = 16383;
defparam ram_block1a84.port_a_logical_ram_depth = 16384;
defparam ram_block1a84.port_a_logical_ram_width = 64;
defparam ram_block1a84.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a84.port_b_address_clear = "none";
defparam ram_block1a84.port_b_address_clock = "clock1";
defparam ram_block1a84.port_b_address_width = 13;
defparam ram_block1a84.port_b_byte_enable_clock = "clock1";
defparam ram_block1a84.port_b_byte_enable_mask_width = 1;
defparam ram_block1a84.port_b_byte_size = 1;
defparam ram_block1a84.port_b_data_in_clock = "clock1";
defparam ram_block1a84.port_b_data_out_clear = "none";
defparam ram_block1a84.port_b_data_out_clock = "none";
defparam ram_block1a84.port_b_data_width = 1;
defparam ram_block1a84.port_b_first_address = 8192;
defparam ram_block1a84.port_b_first_bit_number = 20;
defparam ram_block1a84.port_b_last_address = 16383;
defparam ram_block1a84.port_b_logical_ram_depth = 16384;
defparam ram_block1a84.port_b_logical_ram_width = 64;
defparam ram_block1a84.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a84.port_b_read_enable_clock = "clock1";
defparam ram_block1a84.port_b_write_enable_clock = "clock1";
defparam ram_block1a84.ram_block_type = "auto";
defparam ram_block1a84.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a84.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a84.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a84.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a20(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[20]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus));
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.clk1_core_clock_enable = "ena1";
defparam ram_block1a20.clk1_input_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "bidir_dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 13;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 8191;
defparam ram_block1a20.port_a_logical_ram_depth = 16384;
defparam ram_block1a20.port_a_logical_ram_width = 64;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 13;
defparam ram_block1a20.port_b_byte_enable_clock = "clock1";
defparam ram_block1a20.port_b_byte_enable_mask_width = 1;
defparam ram_block1a20.port_b_byte_size = 1;
defparam ram_block1a20.port_b_data_in_clock = "clock1";
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 8191;
defparam ram_block1a20.port_b_logical_ram_depth = 16384;
defparam ram_block1a20.port_b_logical_ram_width = 64;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.port_b_write_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a20.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a85(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[21]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a85_PORTADATAOUT_bus),
	.portbdataout(ram_block1a85_PORTBDATAOUT_bus));
defparam ram_block1a85.clk0_core_clock_enable = "ena0";
defparam ram_block1a85.clk0_input_clock_enable = "ena0";
defparam ram_block1a85.clk1_core_clock_enable = "ena1";
defparam ram_block1a85.clk1_input_clock_enable = "ena1";
defparam ram_block1a85.data_interleave_offset_in_bits = 1;
defparam ram_block1a85.data_interleave_width_in_bits = 1;
defparam ram_block1a85.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a85.init_file_layout = "port_a";
defparam ram_block1a85.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a85.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a85.operation_mode = "bidir_dual_port";
defparam ram_block1a85.port_a_address_clear = "none";
defparam ram_block1a85.port_a_address_width = 13;
defparam ram_block1a85.port_a_byte_enable_mask_width = 1;
defparam ram_block1a85.port_a_byte_size = 1;
defparam ram_block1a85.port_a_data_out_clear = "none";
defparam ram_block1a85.port_a_data_out_clock = "none";
defparam ram_block1a85.port_a_data_width = 1;
defparam ram_block1a85.port_a_first_address = 8192;
defparam ram_block1a85.port_a_first_bit_number = 21;
defparam ram_block1a85.port_a_last_address = 16383;
defparam ram_block1a85.port_a_logical_ram_depth = 16384;
defparam ram_block1a85.port_a_logical_ram_width = 64;
defparam ram_block1a85.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a85.port_b_address_clear = "none";
defparam ram_block1a85.port_b_address_clock = "clock1";
defparam ram_block1a85.port_b_address_width = 13;
defparam ram_block1a85.port_b_byte_enable_clock = "clock1";
defparam ram_block1a85.port_b_byte_enable_mask_width = 1;
defparam ram_block1a85.port_b_byte_size = 1;
defparam ram_block1a85.port_b_data_in_clock = "clock1";
defparam ram_block1a85.port_b_data_out_clear = "none";
defparam ram_block1a85.port_b_data_out_clock = "none";
defparam ram_block1a85.port_b_data_width = 1;
defparam ram_block1a85.port_b_first_address = 8192;
defparam ram_block1a85.port_b_first_bit_number = 21;
defparam ram_block1a85.port_b_last_address = 16383;
defparam ram_block1a85.port_b_logical_ram_depth = 16384;
defparam ram_block1a85.port_b_logical_ram_width = 64;
defparam ram_block1a85.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a85.port_b_read_enable_clock = "clock1";
defparam ram_block1a85.port_b_write_enable_clock = "clock1";
defparam ram_block1a85.ram_block_type = "auto";
defparam ram_block1a85.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a85.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a85.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a85.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a21(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[21]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus));
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.clk1_core_clock_enable = "ena1";
defparam ram_block1a21.clk1_input_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "bidir_dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 13;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 8191;
defparam ram_block1a21.port_a_logical_ram_depth = 16384;
defparam ram_block1a21.port_a_logical_ram_width = 64;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 13;
defparam ram_block1a21.port_b_byte_enable_clock = "clock1";
defparam ram_block1a21.port_b_byte_enable_mask_width = 1;
defparam ram_block1a21.port_b_byte_size = 1;
defparam ram_block1a21.port_b_data_in_clock = "clock1";
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 8191;
defparam ram_block1a21.port_b_logical_ram_depth = 16384;
defparam ram_block1a21.port_b_logical_ram_width = 64;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.port_b_write_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a21.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a86(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[22]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a86_PORTADATAOUT_bus),
	.portbdataout(ram_block1a86_PORTBDATAOUT_bus));
defparam ram_block1a86.clk0_core_clock_enable = "ena0";
defparam ram_block1a86.clk0_input_clock_enable = "ena0";
defparam ram_block1a86.clk1_core_clock_enable = "ena1";
defparam ram_block1a86.clk1_input_clock_enable = "ena1";
defparam ram_block1a86.data_interleave_offset_in_bits = 1;
defparam ram_block1a86.data_interleave_width_in_bits = 1;
defparam ram_block1a86.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a86.init_file_layout = "port_a";
defparam ram_block1a86.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a86.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a86.operation_mode = "bidir_dual_port";
defparam ram_block1a86.port_a_address_clear = "none";
defparam ram_block1a86.port_a_address_width = 13;
defparam ram_block1a86.port_a_byte_enable_mask_width = 1;
defparam ram_block1a86.port_a_byte_size = 1;
defparam ram_block1a86.port_a_data_out_clear = "none";
defparam ram_block1a86.port_a_data_out_clock = "none";
defparam ram_block1a86.port_a_data_width = 1;
defparam ram_block1a86.port_a_first_address = 8192;
defparam ram_block1a86.port_a_first_bit_number = 22;
defparam ram_block1a86.port_a_last_address = 16383;
defparam ram_block1a86.port_a_logical_ram_depth = 16384;
defparam ram_block1a86.port_a_logical_ram_width = 64;
defparam ram_block1a86.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a86.port_b_address_clear = "none";
defparam ram_block1a86.port_b_address_clock = "clock1";
defparam ram_block1a86.port_b_address_width = 13;
defparam ram_block1a86.port_b_byte_enable_clock = "clock1";
defparam ram_block1a86.port_b_byte_enable_mask_width = 1;
defparam ram_block1a86.port_b_byte_size = 1;
defparam ram_block1a86.port_b_data_in_clock = "clock1";
defparam ram_block1a86.port_b_data_out_clear = "none";
defparam ram_block1a86.port_b_data_out_clock = "none";
defparam ram_block1a86.port_b_data_width = 1;
defparam ram_block1a86.port_b_first_address = 8192;
defparam ram_block1a86.port_b_first_bit_number = 22;
defparam ram_block1a86.port_b_last_address = 16383;
defparam ram_block1a86.port_b_logical_ram_depth = 16384;
defparam ram_block1a86.port_b_logical_ram_width = 64;
defparam ram_block1a86.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a86.port_b_read_enable_clock = "clock1";
defparam ram_block1a86.port_b_write_enable_clock = "clock1";
defparam ram_block1a86.ram_block_type = "auto";
defparam ram_block1a86.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a86.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a86.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a86.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a22(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[22]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus));
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.clk1_core_clock_enable = "ena1";
defparam ram_block1a22.clk1_input_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "bidir_dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 13;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 8191;
defparam ram_block1a22.port_a_logical_ram_depth = 16384;
defparam ram_block1a22.port_a_logical_ram_width = 64;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 13;
defparam ram_block1a22.port_b_byte_enable_clock = "clock1";
defparam ram_block1a22.port_b_byte_enable_mask_width = 1;
defparam ram_block1a22.port_b_byte_size = 1;
defparam ram_block1a22.port_b_data_in_clock = "clock1";
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 8191;
defparam ram_block1a22.port_b_logical_ram_depth = 16384;
defparam ram_block1a22.port_b_logical_ram_width = 64;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.port_b_write_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a22.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a87(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[23]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a87_PORTADATAOUT_bus),
	.portbdataout(ram_block1a87_PORTBDATAOUT_bus));
defparam ram_block1a87.clk0_core_clock_enable = "ena0";
defparam ram_block1a87.clk0_input_clock_enable = "ena0";
defparam ram_block1a87.clk1_core_clock_enable = "ena1";
defparam ram_block1a87.clk1_input_clock_enable = "ena1";
defparam ram_block1a87.data_interleave_offset_in_bits = 1;
defparam ram_block1a87.data_interleave_width_in_bits = 1;
defparam ram_block1a87.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a87.init_file_layout = "port_a";
defparam ram_block1a87.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a87.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a87.operation_mode = "bidir_dual_port";
defparam ram_block1a87.port_a_address_clear = "none";
defparam ram_block1a87.port_a_address_width = 13;
defparam ram_block1a87.port_a_byte_enable_mask_width = 1;
defparam ram_block1a87.port_a_byte_size = 1;
defparam ram_block1a87.port_a_data_out_clear = "none";
defparam ram_block1a87.port_a_data_out_clock = "none";
defparam ram_block1a87.port_a_data_width = 1;
defparam ram_block1a87.port_a_first_address = 8192;
defparam ram_block1a87.port_a_first_bit_number = 23;
defparam ram_block1a87.port_a_last_address = 16383;
defparam ram_block1a87.port_a_logical_ram_depth = 16384;
defparam ram_block1a87.port_a_logical_ram_width = 64;
defparam ram_block1a87.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a87.port_b_address_clear = "none";
defparam ram_block1a87.port_b_address_clock = "clock1";
defparam ram_block1a87.port_b_address_width = 13;
defparam ram_block1a87.port_b_byte_enable_clock = "clock1";
defparam ram_block1a87.port_b_byte_enable_mask_width = 1;
defparam ram_block1a87.port_b_byte_size = 1;
defparam ram_block1a87.port_b_data_in_clock = "clock1";
defparam ram_block1a87.port_b_data_out_clear = "none";
defparam ram_block1a87.port_b_data_out_clock = "none";
defparam ram_block1a87.port_b_data_width = 1;
defparam ram_block1a87.port_b_first_address = 8192;
defparam ram_block1a87.port_b_first_bit_number = 23;
defparam ram_block1a87.port_b_last_address = 16383;
defparam ram_block1a87.port_b_logical_ram_depth = 16384;
defparam ram_block1a87.port_b_logical_ram_width = 64;
defparam ram_block1a87.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a87.port_b_read_enable_clock = "clock1";
defparam ram_block1a87.port_b_write_enable_clock = "clock1";
defparam ram_block1a87.ram_block_type = "auto";
defparam ram_block1a87.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a87.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a87.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a87.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a23(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[23]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[2]}),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus));
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.clk1_core_clock_enable = "ena1";
defparam ram_block1a23.clk1_input_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "bidir_dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 13;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 8191;
defparam ram_block1a23.port_a_logical_ram_depth = 16384;
defparam ram_block1a23.port_a_logical_ram_width = 64;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 13;
defparam ram_block1a23.port_b_byte_enable_clock = "clock1";
defparam ram_block1a23.port_b_byte_enable_mask_width = 1;
defparam ram_block1a23.port_b_byte_size = 1;
defparam ram_block1a23.port_b_data_in_clock = "clock1";
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 8191;
defparam ram_block1a23.port_b_logical_ram_depth = 16384;
defparam ram_block1a23.port_b_logical_ram_width = 64;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.port_b_write_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a23.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a88(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[24]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a88_PORTADATAOUT_bus),
	.portbdataout(ram_block1a88_PORTBDATAOUT_bus));
defparam ram_block1a88.clk0_core_clock_enable = "ena0";
defparam ram_block1a88.clk0_input_clock_enable = "ena0";
defparam ram_block1a88.clk1_core_clock_enable = "ena1";
defparam ram_block1a88.clk1_input_clock_enable = "ena1";
defparam ram_block1a88.data_interleave_offset_in_bits = 1;
defparam ram_block1a88.data_interleave_width_in_bits = 1;
defparam ram_block1a88.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a88.init_file_layout = "port_a";
defparam ram_block1a88.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a88.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a88.operation_mode = "bidir_dual_port";
defparam ram_block1a88.port_a_address_clear = "none";
defparam ram_block1a88.port_a_address_width = 13;
defparam ram_block1a88.port_a_byte_enable_mask_width = 1;
defparam ram_block1a88.port_a_byte_size = 1;
defparam ram_block1a88.port_a_data_out_clear = "none";
defparam ram_block1a88.port_a_data_out_clock = "none";
defparam ram_block1a88.port_a_data_width = 1;
defparam ram_block1a88.port_a_first_address = 8192;
defparam ram_block1a88.port_a_first_bit_number = 24;
defparam ram_block1a88.port_a_last_address = 16383;
defparam ram_block1a88.port_a_logical_ram_depth = 16384;
defparam ram_block1a88.port_a_logical_ram_width = 64;
defparam ram_block1a88.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a88.port_b_address_clear = "none";
defparam ram_block1a88.port_b_address_clock = "clock1";
defparam ram_block1a88.port_b_address_width = 13;
defparam ram_block1a88.port_b_byte_enable_clock = "clock1";
defparam ram_block1a88.port_b_byte_enable_mask_width = 1;
defparam ram_block1a88.port_b_byte_size = 1;
defparam ram_block1a88.port_b_data_in_clock = "clock1";
defparam ram_block1a88.port_b_data_out_clear = "none";
defparam ram_block1a88.port_b_data_out_clock = "none";
defparam ram_block1a88.port_b_data_width = 1;
defparam ram_block1a88.port_b_first_address = 8192;
defparam ram_block1a88.port_b_first_bit_number = 24;
defparam ram_block1a88.port_b_last_address = 16383;
defparam ram_block1a88.port_b_logical_ram_depth = 16384;
defparam ram_block1a88.port_b_logical_ram_width = 64;
defparam ram_block1a88.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a88.port_b_read_enable_clock = "clock1";
defparam ram_block1a88.port_b_write_enable_clock = "clock1";
defparam ram_block1a88.ram_block_type = "auto";
defparam ram_block1a88.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a88.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a88.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a88.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a24(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[24]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus));
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.clk1_core_clock_enable = "ena1";
defparam ram_block1a24.clk1_input_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "bidir_dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 13;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 8191;
defparam ram_block1a24.port_a_logical_ram_depth = 16384;
defparam ram_block1a24.port_a_logical_ram_width = 64;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 13;
defparam ram_block1a24.port_b_byte_enable_clock = "clock1";
defparam ram_block1a24.port_b_byte_enable_mask_width = 1;
defparam ram_block1a24.port_b_byte_size = 1;
defparam ram_block1a24.port_b_data_in_clock = "clock1";
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 8191;
defparam ram_block1a24.port_b_logical_ram_depth = 16384;
defparam ram_block1a24.port_b_logical_ram_width = 64;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.port_b_write_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a89(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[25]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a89_PORTADATAOUT_bus),
	.portbdataout(ram_block1a89_PORTBDATAOUT_bus));
defparam ram_block1a89.clk0_core_clock_enable = "ena0";
defparam ram_block1a89.clk0_input_clock_enable = "ena0";
defparam ram_block1a89.clk1_core_clock_enable = "ena1";
defparam ram_block1a89.clk1_input_clock_enable = "ena1";
defparam ram_block1a89.data_interleave_offset_in_bits = 1;
defparam ram_block1a89.data_interleave_width_in_bits = 1;
defparam ram_block1a89.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a89.init_file_layout = "port_a";
defparam ram_block1a89.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a89.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a89.operation_mode = "bidir_dual_port";
defparam ram_block1a89.port_a_address_clear = "none";
defparam ram_block1a89.port_a_address_width = 13;
defparam ram_block1a89.port_a_byte_enable_mask_width = 1;
defparam ram_block1a89.port_a_byte_size = 1;
defparam ram_block1a89.port_a_data_out_clear = "none";
defparam ram_block1a89.port_a_data_out_clock = "none";
defparam ram_block1a89.port_a_data_width = 1;
defparam ram_block1a89.port_a_first_address = 8192;
defparam ram_block1a89.port_a_first_bit_number = 25;
defparam ram_block1a89.port_a_last_address = 16383;
defparam ram_block1a89.port_a_logical_ram_depth = 16384;
defparam ram_block1a89.port_a_logical_ram_width = 64;
defparam ram_block1a89.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a89.port_b_address_clear = "none";
defparam ram_block1a89.port_b_address_clock = "clock1";
defparam ram_block1a89.port_b_address_width = 13;
defparam ram_block1a89.port_b_byte_enable_clock = "clock1";
defparam ram_block1a89.port_b_byte_enable_mask_width = 1;
defparam ram_block1a89.port_b_byte_size = 1;
defparam ram_block1a89.port_b_data_in_clock = "clock1";
defparam ram_block1a89.port_b_data_out_clear = "none";
defparam ram_block1a89.port_b_data_out_clock = "none";
defparam ram_block1a89.port_b_data_width = 1;
defparam ram_block1a89.port_b_first_address = 8192;
defparam ram_block1a89.port_b_first_bit_number = 25;
defparam ram_block1a89.port_b_last_address = 16383;
defparam ram_block1a89.port_b_logical_ram_depth = 16384;
defparam ram_block1a89.port_b_logical_ram_width = 64;
defparam ram_block1a89.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a89.port_b_read_enable_clock = "clock1";
defparam ram_block1a89.port_b_write_enable_clock = "clock1";
defparam ram_block1a89.ram_block_type = "auto";
defparam ram_block1a89.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a89.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a89.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a89.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a25(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[25]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus));
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.clk1_core_clock_enable = "ena1";
defparam ram_block1a25.clk1_input_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "bidir_dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 13;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 8191;
defparam ram_block1a25.port_a_logical_ram_depth = 16384;
defparam ram_block1a25.port_a_logical_ram_width = 64;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 13;
defparam ram_block1a25.port_b_byte_enable_clock = "clock1";
defparam ram_block1a25.port_b_byte_enable_mask_width = 1;
defparam ram_block1a25.port_b_byte_size = 1;
defparam ram_block1a25.port_b_data_in_clock = "clock1";
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 8191;
defparam ram_block1a25.port_b_logical_ram_depth = 16384;
defparam ram_block1a25.port_b_logical_ram_width = 64;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.port_b_write_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a25.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a90(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[26]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a90_PORTADATAOUT_bus),
	.portbdataout(ram_block1a90_PORTBDATAOUT_bus));
defparam ram_block1a90.clk0_core_clock_enable = "ena0";
defparam ram_block1a90.clk0_input_clock_enable = "ena0";
defparam ram_block1a90.clk1_core_clock_enable = "ena1";
defparam ram_block1a90.clk1_input_clock_enable = "ena1";
defparam ram_block1a90.data_interleave_offset_in_bits = 1;
defparam ram_block1a90.data_interleave_width_in_bits = 1;
defparam ram_block1a90.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a90.init_file_layout = "port_a";
defparam ram_block1a90.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a90.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a90.operation_mode = "bidir_dual_port";
defparam ram_block1a90.port_a_address_clear = "none";
defparam ram_block1a90.port_a_address_width = 13;
defparam ram_block1a90.port_a_byte_enable_mask_width = 1;
defparam ram_block1a90.port_a_byte_size = 1;
defparam ram_block1a90.port_a_data_out_clear = "none";
defparam ram_block1a90.port_a_data_out_clock = "none";
defparam ram_block1a90.port_a_data_width = 1;
defparam ram_block1a90.port_a_first_address = 8192;
defparam ram_block1a90.port_a_first_bit_number = 26;
defparam ram_block1a90.port_a_last_address = 16383;
defparam ram_block1a90.port_a_logical_ram_depth = 16384;
defparam ram_block1a90.port_a_logical_ram_width = 64;
defparam ram_block1a90.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a90.port_b_address_clear = "none";
defparam ram_block1a90.port_b_address_clock = "clock1";
defparam ram_block1a90.port_b_address_width = 13;
defparam ram_block1a90.port_b_byte_enable_clock = "clock1";
defparam ram_block1a90.port_b_byte_enable_mask_width = 1;
defparam ram_block1a90.port_b_byte_size = 1;
defparam ram_block1a90.port_b_data_in_clock = "clock1";
defparam ram_block1a90.port_b_data_out_clear = "none";
defparam ram_block1a90.port_b_data_out_clock = "none";
defparam ram_block1a90.port_b_data_width = 1;
defparam ram_block1a90.port_b_first_address = 8192;
defparam ram_block1a90.port_b_first_bit_number = 26;
defparam ram_block1a90.port_b_last_address = 16383;
defparam ram_block1a90.port_b_logical_ram_depth = 16384;
defparam ram_block1a90.port_b_logical_ram_width = 64;
defparam ram_block1a90.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a90.port_b_read_enable_clock = "clock1";
defparam ram_block1a90.port_b_write_enable_clock = "clock1";
defparam ram_block1a90.ram_block_type = "auto";
defparam ram_block1a90.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a90.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a90.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a90.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a26(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[26]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus));
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.clk1_core_clock_enable = "ena1";
defparam ram_block1a26.clk1_input_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "bidir_dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 13;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 8191;
defparam ram_block1a26.port_a_logical_ram_depth = 16384;
defparam ram_block1a26.port_a_logical_ram_width = 64;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 13;
defparam ram_block1a26.port_b_byte_enable_clock = "clock1";
defparam ram_block1a26.port_b_byte_enable_mask_width = 1;
defparam ram_block1a26.port_b_byte_size = 1;
defparam ram_block1a26.port_b_data_in_clock = "clock1";
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 8191;
defparam ram_block1a26.port_b_logical_ram_depth = 16384;
defparam ram_block1a26.port_b_logical_ram_width = 64;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.port_b_write_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a91(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[27]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a91_PORTADATAOUT_bus),
	.portbdataout(ram_block1a91_PORTBDATAOUT_bus));
defparam ram_block1a91.clk0_core_clock_enable = "ena0";
defparam ram_block1a91.clk0_input_clock_enable = "ena0";
defparam ram_block1a91.clk1_core_clock_enable = "ena1";
defparam ram_block1a91.clk1_input_clock_enable = "ena1";
defparam ram_block1a91.data_interleave_offset_in_bits = 1;
defparam ram_block1a91.data_interleave_width_in_bits = 1;
defparam ram_block1a91.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a91.init_file_layout = "port_a";
defparam ram_block1a91.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a91.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a91.operation_mode = "bidir_dual_port";
defparam ram_block1a91.port_a_address_clear = "none";
defparam ram_block1a91.port_a_address_width = 13;
defparam ram_block1a91.port_a_byte_enable_mask_width = 1;
defparam ram_block1a91.port_a_byte_size = 1;
defparam ram_block1a91.port_a_data_out_clear = "none";
defparam ram_block1a91.port_a_data_out_clock = "none";
defparam ram_block1a91.port_a_data_width = 1;
defparam ram_block1a91.port_a_first_address = 8192;
defparam ram_block1a91.port_a_first_bit_number = 27;
defparam ram_block1a91.port_a_last_address = 16383;
defparam ram_block1a91.port_a_logical_ram_depth = 16384;
defparam ram_block1a91.port_a_logical_ram_width = 64;
defparam ram_block1a91.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a91.port_b_address_clear = "none";
defparam ram_block1a91.port_b_address_clock = "clock1";
defparam ram_block1a91.port_b_address_width = 13;
defparam ram_block1a91.port_b_byte_enable_clock = "clock1";
defparam ram_block1a91.port_b_byte_enable_mask_width = 1;
defparam ram_block1a91.port_b_byte_size = 1;
defparam ram_block1a91.port_b_data_in_clock = "clock1";
defparam ram_block1a91.port_b_data_out_clear = "none";
defparam ram_block1a91.port_b_data_out_clock = "none";
defparam ram_block1a91.port_b_data_width = 1;
defparam ram_block1a91.port_b_first_address = 8192;
defparam ram_block1a91.port_b_first_bit_number = 27;
defparam ram_block1a91.port_b_last_address = 16383;
defparam ram_block1a91.port_b_logical_ram_depth = 16384;
defparam ram_block1a91.port_b_logical_ram_width = 64;
defparam ram_block1a91.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a91.port_b_read_enable_clock = "clock1";
defparam ram_block1a91.port_b_write_enable_clock = "clock1";
defparam ram_block1a91.ram_block_type = "auto";
defparam ram_block1a91.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a91.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a91.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a91.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a27(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[27]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus));
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.clk1_core_clock_enable = "ena1";
defparam ram_block1a27.clk1_input_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "bidir_dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 13;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 8191;
defparam ram_block1a27.port_a_logical_ram_depth = 16384;
defparam ram_block1a27.port_a_logical_ram_width = 64;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 13;
defparam ram_block1a27.port_b_byte_enable_clock = "clock1";
defparam ram_block1a27.port_b_byte_enable_mask_width = 1;
defparam ram_block1a27.port_b_byte_size = 1;
defparam ram_block1a27.port_b_data_in_clock = "clock1";
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 8191;
defparam ram_block1a27.port_b_logical_ram_depth = 16384;
defparam ram_block1a27.port_b_logical_ram_width = 64;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.port_b_write_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a27.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a92(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[28]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a92_PORTADATAOUT_bus),
	.portbdataout(ram_block1a92_PORTBDATAOUT_bus));
defparam ram_block1a92.clk0_core_clock_enable = "ena0";
defparam ram_block1a92.clk0_input_clock_enable = "ena0";
defparam ram_block1a92.clk1_core_clock_enable = "ena1";
defparam ram_block1a92.clk1_input_clock_enable = "ena1";
defparam ram_block1a92.data_interleave_offset_in_bits = 1;
defparam ram_block1a92.data_interleave_width_in_bits = 1;
defparam ram_block1a92.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a92.init_file_layout = "port_a";
defparam ram_block1a92.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a92.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a92.operation_mode = "bidir_dual_port";
defparam ram_block1a92.port_a_address_clear = "none";
defparam ram_block1a92.port_a_address_width = 13;
defparam ram_block1a92.port_a_byte_enable_mask_width = 1;
defparam ram_block1a92.port_a_byte_size = 1;
defparam ram_block1a92.port_a_data_out_clear = "none";
defparam ram_block1a92.port_a_data_out_clock = "none";
defparam ram_block1a92.port_a_data_width = 1;
defparam ram_block1a92.port_a_first_address = 8192;
defparam ram_block1a92.port_a_first_bit_number = 28;
defparam ram_block1a92.port_a_last_address = 16383;
defparam ram_block1a92.port_a_logical_ram_depth = 16384;
defparam ram_block1a92.port_a_logical_ram_width = 64;
defparam ram_block1a92.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a92.port_b_address_clear = "none";
defparam ram_block1a92.port_b_address_clock = "clock1";
defparam ram_block1a92.port_b_address_width = 13;
defparam ram_block1a92.port_b_byte_enable_clock = "clock1";
defparam ram_block1a92.port_b_byte_enable_mask_width = 1;
defparam ram_block1a92.port_b_byte_size = 1;
defparam ram_block1a92.port_b_data_in_clock = "clock1";
defparam ram_block1a92.port_b_data_out_clear = "none";
defparam ram_block1a92.port_b_data_out_clock = "none";
defparam ram_block1a92.port_b_data_width = 1;
defparam ram_block1a92.port_b_first_address = 8192;
defparam ram_block1a92.port_b_first_bit_number = 28;
defparam ram_block1a92.port_b_last_address = 16383;
defparam ram_block1a92.port_b_logical_ram_depth = 16384;
defparam ram_block1a92.port_b_logical_ram_width = 64;
defparam ram_block1a92.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a92.port_b_read_enable_clock = "clock1";
defparam ram_block1a92.port_b_write_enable_clock = "clock1";
defparam ram_block1a92.ram_block_type = "auto";
defparam ram_block1a92.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a92.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a92.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a92.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a28(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[28]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus));
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.clk1_core_clock_enable = "ena1";
defparam ram_block1a28.clk1_input_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "bidir_dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 13;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 8191;
defparam ram_block1a28.port_a_logical_ram_depth = 16384;
defparam ram_block1a28.port_a_logical_ram_width = 64;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 13;
defparam ram_block1a28.port_b_byte_enable_clock = "clock1";
defparam ram_block1a28.port_b_byte_enable_mask_width = 1;
defparam ram_block1a28.port_b_byte_size = 1;
defparam ram_block1a28.port_b_data_in_clock = "clock1";
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 8191;
defparam ram_block1a28.port_b_logical_ram_depth = 16384;
defparam ram_block1a28.port_b_logical_ram_width = 64;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.port_b_write_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a28.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a93(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[29]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a93_PORTADATAOUT_bus),
	.portbdataout(ram_block1a93_PORTBDATAOUT_bus));
defparam ram_block1a93.clk0_core_clock_enable = "ena0";
defparam ram_block1a93.clk0_input_clock_enable = "ena0";
defparam ram_block1a93.clk1_core_clock_enable = "ena1";
defparam ram_block1a93.clk1_input_clock_enable = "ena1";
defparam ram_block1a93.data_interleave_offset_in_bits = 1;
defparam ram_block1a93.data_interleave_width_in_bits = 1;
defparam ram_block1a93.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a93.init_file_layout = "port_a";
defparam ram_block1a93.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a93.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a93.operation_mode = "bidir_dual_port";
defparam ram_block1a93.port_a_address_clear = "none";
defparam ram_block1a93.port_a_address_width = 13;
defparam ram_block1a93.port_a_byte_enable_mask_width = 1;
defparam ram_block1a93.port_a_byte_size = 1;
defparam ram_block1a93.port_a_data_out_clear = "none";
defparam ram_block1a93.port_a_data_out_clock = "none";
defparam ram_block1a93.port_a_data_width = 1;
defparam ram_block1a93.port_a_first_address = 8192;
defparam ram_block1a93.port_a_first_bit_number = 29;
defparam ram_block1a93.port_a_last_address = 16383;
defparam ram_block1a93.port_a_logical_ram_depth = 16384;
defparam ram_block1a93.port_a_logical_ram_width = 64;
defparam ram_block1a93.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a93.port_b_address_clear = "none";
defparam ram_block1a93.port_b_address_clock = "clock1";
defparam ram_block1a93.port_b_address_width = 13;
defparam ram_block1a93.port_b_byte_enable_clock = "clock1";
defparam ram_block1a93.port_b_byte_enable_mask_width = 1;
defparam ram_block1a93.port_b_byte_size = 1;
defparam ram_block1a93.port_b_data_in_clock = "clock1";
defparam ram_block1a93.port_b_data_out_clear = "none";
defparam ram_block1a93.port_b_data_out_clock = "none";
defparam ram_block1a93.port_b_data_width = 1;
defparam ram_block1a93.port_b_first_address = 8192;
defparam ram_block1a93.port_b_first_bit_number = 29;
defparam ram_block1a93.port_b_last_address = 16383;
defparam ram_block1a93.port_b_logical_ram_depth = 16384;
defparam ram_block1a93.port_b_logical_ram_width = 64;
defparam ram_block1a93.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a93.port_b_read_enable_clock = "clock1";
defparam ram_block1a93.port_b_write_enable_clock = "clock1";
defparam ram_block1a93.ram_block_type = "auto";
defparam ram_block1a93.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a93.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a93.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a93.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a29(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[29]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus));
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.clk1_core_clock_enable = "ena1";
defparam ram_block1a29.clk1_input_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "bidir_dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 13;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 8191;
defparam ram_block1a29.port_a_logical_ram_depth = 16384;
defparam ram_block1a29.port_a_logical_ram_width = 64;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 13;
defparam ram_block1a29.port_b_byte_enable_clock = "clock1";
defparam ram_block1a29.port_b_byte_enable_mask_width = 1;
defparam ram_block1a29.port_b_byte_size = 1;
defparam ram_block1a29.port_b_data_in_clock = "clock1";
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 8191;
defparam ram_block1a29.port_b_logical_ram_depth = 16384;
defparam ram_block1a29.port_b_logical_ram_width = 64;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.port_b_write_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a29.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a94(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[30]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a94_PORTADATAOUT_bus),
	.portbdataout(ram_block1a94_PORTBDATAOUT_bus));
defparam ram_block1a94.clk0_core_clock_enable = "ena0";
defparam ram_block1a94.clk0_input_clock_enable = "ena0";
defparam ram_block1a94.clk1_core_clock_enable = "ena1";
defparam ram_block1a94.clk1_input_clock_enable = "ena1";
defparam ram_block1a94.data_interleave_offset_in_bits = 1;
defparam ram_block1a94.data_interleave_width_in_bits = 1;
defparam ram_block1a94.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a94.init_file_layout = "port_a";
defparam ram_block1a94.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a94.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a94.operation_mode = "bidir_dual_port";
defparam ram_block1a94.port_a_address_clear = "none";
defparam ram_block1a94.port_a_address_width = 13;
defparam ram_block1a94.port_a_byte_enable_mask_width = 1;
defparam ram_block1a94.port_a_byte_size = 1;
defparam ram_block1a94.port_a_data_out_clear = "none";
defparam ram_block1a94.port_a_data_out_clock = "none";
defparam ram_block1a94.port_a_data_width = 1;
defparam ram_block1a94.port_a_first_address = 8192;
defparam ram_block1a94.port_a_first_bit_number = 30;
defparam ram_block1a94.port_a_last_address = 16383;
defparam ram_block1a94.port_a_logical_ram_depth = 16384;
defparam ram_block1a94.port_a_logical_ram_width = 64;
defparam ram_block1a94.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a94.port_b_address_clear = "none";
defparam ram_block1a94.port_b_address_clock = "clock1";
defparam ram_block1a94.port_b_address_width = 13;
defparam ram_block1a94.port_b_byte_enable_clock = "clock1";
defparam ram_block1a94.port_b_byte_enable_mask_width = 1;
defparam ram_block1a94.port_b_byte_size = 1;
defparam ram_block1a94.port_b_data_in_clock = "clock1";
defparam ram_block1a94.port_b_data_out_clear = "none";
defparam ram_block1a94.port_b_data_out_clock = "none";
defparam ram_block1a94.port_b_data_width = 1;
defparam ram_block1a94.port_b_first_address = 8192;
defparam ram_block1a94.port_b_first_bit_number = 30;
defparam ram_block1a94.port_b_last_address = 16383;
defparam ram_block1a94.port_b_logical_ram_depth = 16384;
defparam ram_block1a94.port_b_logical_ram_width = 64;
defparam ram_block1a94.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a94.port_b_read_enable_clock = "clock1";
defparam ram_block1a94.port_b_write_enable_clock = "clock1";
defparam ram_block1a94.ram_block_type = "auto";
defparam ram_block1a94.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a94.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a94.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a94.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a30(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[30]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus));
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.clk1_core_clock_enable = "ena1";
defparam ram_block1a30.clk1_input_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "bidir_dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 13;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 8191;
defparam ram_block1a30.port_a_logical_ram_depth = 16384;
defparam ram_block1a30.port_a_logical_ram_width = 64;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 13;
defparam ram_block1a30.port_b_byte_enable_clock = "clock1";
defparam ram_block1a30.port_b_byte_enable_mask_width = 1;
defparam ram_block1a30.port_b_byte_size = 1;
defparam ram_block1a30.port_b_data_in_clock = "clock1";
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 8191;
defparam ram_block1a30.port_b_logical_ram_depth = 16384;
defparam ram_block1a30.port_b_logical_ram_width = 64;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.port_b_write_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a95(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[31]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a95_PORTADATAOUT_bus),
	.portbdataout(ram_block1a95_PORTBDATAOUT_bus));
defparam ram_block1a95.clk0_core_clock_enable = "ena0";
defparam ram_block1a95.clk0_input_clock_enable = "ena0";
defparam ram_block1a95.clk1_core_clock_enable = "ena1";
defparam ram_block1a95.clk1_input_clock_enable = "ena1";
defparam ram_block1a95.data_interleave_offset_in_bits = 1;
defparam ram_block1a95.data_interleave_width_in_bits = 1;
defparam ram_block1a95.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a95.init_file_layout = "port_a";
defparam ram_block1a95.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a95.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a95.operation_mode = "bidir_dual_port";
defparam ram_block1a95.port_a_address_clear = "none";
defparam ram_block1a95.port_a_address_width = 13;
defparam ram_block1a95.port_a_byte_enable_mask_width = 1;
defparam ram_block1a95.port_a_byte_size = 1;
defparam ram_block1a95.port_a_data_out_clear = "none";
defparam ram_block1a95.port_a_data_out_clock = "none";
defparam ram_block1a95.port_a_data_width = 1;
defparam ram_block1a95.port_a_first_address = 8192;
defparam ram_block1a95.port_a_first_bit_number = 31;
defparam ram_block1a95.port_a_last_address = 16383;
defparam ram_block1a95.port_a_logical_ram_depth = 16384;
defparam ram_block1a95.port_a_logical_ram_width = 64;
defparam ram_block1a95.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a95.port_b_address_clear = "none";
defparam ram_block1a95.port_b_address_clock = "clock1";
defparam ram_block1a95.port_b_address_width = 13;
defparam ram_block1a95.port_b_byte_enable_clock = "clock1";
defparam ram_block1a95.port_b_byte_enable_mask_width = 1;
defparam ram_block1a95.port_b_byte_size = 1;
defparam ram_block1a95.port_b_data_in_clock = "clock1";
defparam ram_block1a95.port_b_data_out_clear = "none";
defparam ram_block1a95.port_b_data_out_clock = "none";
defparam ram_block1a95.port_b_data_width = 1;
defparam ram_block1a95.port_b_first_address = 8192;
defparam ram_block1a95.port_b_first_bit_number = 31;
defparam ram_block1a95.port_b_last_address = 16383;
defparam ram_block1a95.port_b_logical_ram_depth = 16384;
defparam ram_block1a95.port_b_logical_ram_width = 64;
defparam ram_block1a95.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a95.port_b_read_enable_clock = "clock1";
defparam ram_block1a95.port_b_write_enable_clock = "clock1";
defparam ram_block1a95.ram_block_type = "auto";
defparam ram_block1a95.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a95.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a95.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a95.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a31(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[31]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[3]}),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus));
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.clk1_core_clock_enable = "ena1";
defparam ram_block1a31.clk1_input_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "bidir_dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 13;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 8191;
defparam ram_block1a31.port_a_logical_ram_depth = 16384;
defparam ram_block1a31.port_a_logical_ram_width = 64;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 13;
defparam ram_block1a31.port_b_byte_enable_clock = "clock1";
defparam ram_block1a31.port_b_byte_enable_mask_width = 1;
defparam ram_block1a31.port_b_byte_size = 1;
defparam ram_block1a31.port_b_data_in_clock = "clock1";
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 8191;
defparam ram_block1a31.port_b_logical_ram_depth = 16384;
defparam ram_block1a31.port_b_logical_ram_width = 64;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.port_b_write_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a31.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a96(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[32]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[32]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a96_PORTADATAOUT_bus),
	.portbdataout(ram_block1a96_PORTBDATAOUT_bus));
defparam ram_block1a96.clk0_core_clock_enable = "ena0";
defparam ram_block1a96.clk0_input_clock_enable = "ena0";
defparam ram_block1a96.clk1_core_clock_enable = "ena1";
defparam ram_block1a96.clk1_input_clock_enable = "ena1";
defparam ram_block1a96.data_interleave_offset_in_bits = 1;
defparam ram_block1a96.data_interleave_width_in_bits = 1;
defparam ram_block1a96.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a96.init_file_layout = "port_a";
defparam ram_block1a96.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a96.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a96.operation_mode = "bidir_dual_port";
defparam ram_block1a96.port_a_address_clear = "none";
defparam ram_block1a96.port_a_address_width = 13;
defparam ram_block1a96.port_a_byte_enable_mask_width = 1;
defparam ram_block1a96.port_a_byte_size = 1;
defparam ram_block1a96.port_a_data_out_clear = "none";
defparam ram_block1a96.port_a_data_out_clock = "none";
defparam ram_block1a96.port_a_data_width = 1;
defparam ram_block1a96.port_a_first_address = 8192;
defparam ram_block1a96.port_a_first_bit_number = 32;
defparam ram_block1a96.port_a_last_address = 16383;
defparam ram_block1a96.port_a_logical_ram_depth = 16384;
defparam ram_block1a96.port_a_logical_ram_width = 64;
defparam ram_block1a96.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a96.port_b_address_clear = "none";
defparam ram_block1a96.port_b_address_clock = "clock1";
defparam ram_block1a96.port_b_address_width = 13;
defparam ram_block1a96.port_b_byte_enable_clock = "clock1";
defparam ram_block1a96.port_b_byte_enable_mask_width = 1;
defparam ram_block1a96.port_b_byte_size = 1;
defparam ram_block1a96.port_b_data_in_clock = "clock1";
defparam ram_block1a96.port_b_data_out_clear = "none";
defparam ram_block1a96.port_b_data_out_clock = "none";
defparam ram_block1a96.port_b_data_width = 1;
defparam ram_block1a96.port_b_first_address = 8192;
defparam ram_block1a96.port_b_first_bit_number = 32;
defparam ram_block1a96.port_b_last_address = 16383;
defparam ram_block1a96.port_b_logical_ram_depth = 16384;
defparam ram_block1a96.port_b_logical_ram_width = 64;
defparam ram_block1a96.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a96.port_b_read_enable_clock = "clock1";
defparam ram_block1a96.port_b_write_enable_clock = "clock1";
defparam ram_block1a96.ram_block_type = "auto";
defparam ram_block1a96.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a96.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a96.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a96.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a32(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[32]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[32]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a32_PORTADATAOUT_bus),
	.portbdataout(ram_block1a32_PORTBDATAOUT_bus));
defparam ram_block1a32.clk0_core_clock_enable = "ena0";
defparam ram_block1a32.clk0_input_clock_enable = "ena0";
defparam ram_block1a32.clk1_core_clock_enable = "ena1";
defparam ram_block1a32.clk1_input_clock_enable = "ena1";
defparam ram_block1a32.data_interleave_offset_in_bits = 1;
defparam ram_block1a32.data_interleave_width_in_bits = 1;
defparam ram_block1a32.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a32.init_file_layout = "port_a";
defparam ram_block1a32.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a32.operation_mode = "bidir_dual_port";
defparam ram_block1a32.port_a_address_clear = "none";
defparam ram_block1a32.port_a_address_width = 13;
defparam ram_block1a32.port_a_byte_enable_mask_width = 1;
defparam ram_block1a32.port_a_byte_size = 1;
defparam ram_block1a32.port_a_data_out_clear = "none";
defparam ram_block1a32.port_a_data_out_clock = "none";
defparam ram_block1a32.port_a_data_width = 1;
defparam ram_block1a32.port_a_first_address = 0;
defparam ram_block1a32.port_a_first_bit_number = 32;
defparam ram_block1a32.port_a_last_address = 8191;
defparam ram_block1a32.port_a_logical_ram_depth = 16384;
defparam ram_block1a32.port_a_logical_ram_width = 64;
defparam ram_block1a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a32.port_b_address_clear = "none";
defparam ram_block1a32.port_b_address_clock = "clock1";
defparam ram_block1a32.port_b_address_width = 13;
defparam ram_block1a32.port_b_byte_enable_clock = "clock1";
defparam ram_block1a32.port_b_byte_enable_mask_width = 1;
defparam ram_block1a32.port_b_byte_size = 1;
defparam ram_block1a32.port_b_data_in_clock = "clock1";
defparam ram_block1a32.port_b_data_out_clear = "none";
defparam ram_block1a32.port_b_data_out_clock = "none";
defparam ram_block1a32.port_b_data_width = 1;
defparam ram_block1a32.port_b_first_address = 0;
defparam ram_block1a32.port_b_first_bit_number = 32;
defparam ram_block1a32.port_b_last_address = 8191;
defparam ram_block1a32.port_b_logical_ram_depth = 16384;
defparam ram_block1a32.port_b_logical_ram_width = 64;
defparam ram_block1a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a32.port_b_read_enable_clock = "clock1";
defparam ram_block1a32.port_b_write_enable_clock = "clock1";
defparam ram_block1a32.ram_block_type = "auto";
defparam ram_block1a32.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a32.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a32.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a32.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a97(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[33]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[33]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a97_PORTADATAOUT_bus),
	.portbdataout(ram_block1a97_PORTBDATAOUT_bus));
defparam ram_block1a97.clk0_core_clock_enable = "ena0";
defparam ram_block1a97.clk0_input_clock_enable = "ena0";
defparam ram_block1a97.clk1_core_clock_enable = "ena1";
defparam ram_block1a97.clk1_input_clock_enable = "ena1";
defparam ram_block1a97.data_interleave_offset_in_bits = 1;
defparam ram_block1a97.data_interleave_width_in_bits = 1;
defparam ram_block1a97.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a97.init_file_layout = "port_a";
defparam ram_block1a97.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a97.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a97.operation_mode = "bidir_dual_port";
defparam ram_block1a97.port_a_address_clear = "none";
defparam ram_block1a97.port_a_address_width = 13;
defparam ram_block1a97.port_a_byte_enable_mask_width = 1;
defparam ram_block1a97.port_a_byte_size = 1;
defparam ram_block1a97.port_a_data_out_clear = "none";
defparam ram_block1a97.port_a_data_out_clock = "none";
defparam ram_block1a97.port_a_data_width = 1;
defparam ram_block1a97.port_a_first_address = 8192;
defparam ram_block1a97.port_a_first_bit_number = 33;
defparam ram_block1a97.port_a_last_address = 16383;
defparam ram_block1a97.port_a_logical_ram_depth = 16384;
defparam ram_block1a97.port_a_logical_ram_width = 64;
defparam ram_block1a97.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a97.port_b_address_clear = "none";
defparam ram_block1a97.port_b_address_clock = "clock1";
defparam ram_block1a97.port_b_address_width = 13;
defparam ram_block1a97.port_b_byte_enable_clock = "clock1";
defparam ram_block1a97.port_b_byte_enable_mask_width = 1;
defparam ram_block1a97.port_b_byte_size = 1;
defparam ram_block1a97.port_b_data_in_clock = "clock1";
defparam ram_block1a97.port_b_data_out_clear = "none";
defparam ram_block1a97.port_b_data_out_clock = "none";
defparam ram_block1a97.port_b_data_width = 1;
defparam ram_block1a97.port_b_first_address = 8192;
defparam ram_block1a97.port_b_first_bit_number = 33;
defparam ram_block1a97.port_b_last_address = 16383;
defparam ram_block1a97.port_b_logical_ram_depth = 16384;
defparam ram_block1a97.port_b_logical_ram_width = 64;
defparam ram_block1a97.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a97.port_b_read_enable_clock = "clock1";
defparam ram_block1a97.port_b_write_enable_clock = "clock1";
defparam ram_block1a97.ram_block_type = "auto";
defparam ram_block1a97.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a97.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a97.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a97.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a33(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[33]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[33]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a33_PORTADATAOUT_bus),
	.portbdataout(ram_block1a33_PORTBDATAOUT_bus));
defparam ram_block1a33.clk0_core_clock_enable = "ena0";
defparam ram_block1a33.clk0_input_clock_enable = "ena0";
defparam ram_block1a33.clk1_core_clock_enable = "ena1";
defparam ram_block1a33.clk1_input_clock_enable = "ena1";
defparam ram_block1a33.data_interleave_offset_in_bits = 1;
defparam ram_block1a33.data_interleave_width_in_bits = 1;
defparam ram_block1a33.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a33.init_file_layout = "port_a";
defparam ram_block1a33.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a33.operation_mode = "bidir_dual_port";
defparam ram_block1a33.port_a_address_clear = "none";
defparam ram_block1a33.port_a_address_width = 13;
defparam ram_block1a33.port_a_byte_enable_mask_width = 1;
defparam ram_block1a33.port_a_byte_size = 1;
defparam ram_block1a33.port_a_data_out_clear = "none";
defparam ram_block1a33.port_a_data_out_clock = "none";
defparam ram_block1a33.port_a_data_width = 1;
defparam ram_block1a33.port_a_first_address = 0;
defparam ram_block1a33.port_a_first_bit_number = 33;
defparam ram_block1a33.port_a_last_address = 8191;
defparam ram_block1a33.port_a_logical_ram_depth = 16384;
defparam ram_block1a33.port_a_logical_ram_width = 64;
defparam ram_block1a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a33.port_b_address_clear = "none";
defparam ram_block1a33.port_b_address_clock = "clock1";
defparam ram_block1a33.port_b_address_width = 13;
defparam ram_block1a33.port_b_byte_enable_clock = "clock1";
defparam ram_block1a33.port_b_byte_enable_mask_width = 1;
defparam ram_block1a33.port_b_byte_size = 1;
defparam ram_block1a33.port_b_data_in_clock = "clock1";
defparam ram_block1a33.port_b_data_out_clear = "none";
defparam ram_block1a33.port_b_data_out_clock = "none";
defparam ram_block1a33.port_b_data_width = 1;
defparam ram_block1a33.port_b_first_address = 0;
defparam ram_block1a33.port_b_first_bit_number = 33;
defparam ram_block1a33.port_b_last_address = 8191;
defparam ram_block1a33.port_b_logical_ram_depth = 16384;
defparam ram_block1a33.port_b_logical_ram_width = 64;
defparam ram_block1a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a33.port_b_read_enable_clock = "clock1";
defparam ram_block1a33.port_b_write_enable_clock = "clock1";
defparam ram_block1a33.ram_block_type = "auto";
defparam ram_block1a33.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a33.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a33.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a33.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a98(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[34]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[34]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a98_PORTADATAOUT_bus),
	.portbdataout(ram_block1a98_PORTBDATAOUT_bus));
defparam ram_block1a98.clk0_core_clock_enable = "ena0";
defparam ram_block1a98.clk0_input_clock_enable = "ena0";
defparam ram_block1a98.clk1_core_clock_enable = "ena1";
defparam ram_block1a98.clk1_input_clock_enable = "ena1";
defparam ram_block1a98.data_interleave_offset_in_bits = 1;
defparam ram_block1a98.data_interleave_width_in_bits = 1;
defparam ram_block1a98.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a98.init_file_layout = "port_a";
defparam ram_block1a98.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a98.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a98.operation_mode = "bidir_dual_port";
defparam ram_block1a98.port_a_address_clear = "none";
defparam ram_block1a98.port_a_address_width = 13;
defparam ram_block1a98.port_a_byte_enable_mask_width = 1;
defparam ram_block1a98.port_a_byte_size = 1;
defparam ram_block1a98.port_a_data_out_clear = "none";
defparam ram_block1a98.port_a_data_out_clock = "none";
defparam ram_block1a98.port_a_data_width = 1;
defparam ram_block1a98.port_a_first_address = 8192;
defparam ram_block1a98.port_a_first_bit_number = 34;
defparam ram_block1a98.port_a_last_address = 16383;
defparam ram_block1a98.port_a_logical_ram_depth = 16384;
defparam ram_block1a98.port_a_logical_ram_width = 64;
defparam ram_block1a98.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a98.port_b_address_clear = "none";
defparam ram_block1a98.port_b_address_clock = "clock1";
defparam ram_block1a98.port_b_address_width = 13;
defparam ram_block1a98.port_b_byte_enable_clock = "clock1";
defparam ram_block1a98.port_b_byte_enable_mask_width = 1;
defparam ram_block1a98.port_b_byte_size = 1;
defparam ram_block1a98.port_b_data_in_clock = "clock1";
defparam ram_block1a98.port_b_data_out_clear = "none";
defparam ram_block1a98.port_b_data_out_clock = "none";
defparam ram_block1a98.port_b_data_width = 1;
defparam ram_block1a98.port_b_first_address = 8192;
defparam ram_block1a98.port_b_first_bit_number = 34;
defparam ram_block1a98.port_b_last_address = 16383;
defparam ram_block1a98.port_b_logical_ram_depth = 16384;
defparam ram_block1a98.port_b_logical_ram_width = 64;
defparam ram_block1a98.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a98.port_b_read_enable_clock = "clock1";
defparam ram_block1a98.port_b_write_enable_clock = "clock1";
defparam ram_block1a98.ram_block_type = "auto";
defparam ram_block1a98.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a98.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a98.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a98.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a34(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[34]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[34]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a34_PORTADATAOUT_bus),
	.portbdataout(ram_block1a34_PORTBDATAOUT_bus));
defparam ram_block1a34.clk0_core_clock_enable = "ena0";
defparam ram_block1a34.clk0_input_clock_enable = "ena0";
defparam ram_block1a34.clk1_core_clock_enable = "ena1";
defparam ram_block1a34.clk1_input_clock_enable = "ena1";
defparam ram_block1a34.data_interleave_offset_in_bits = 1;
defparam ram_block1a34.data_interleave_width_in_bits = 1;
defparam ram_block1a34.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a34.init_file_layout = "port_a";
defparam ram_block1a34.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a34.operation_mode = "bidir_dual_port";
defparam ram_block1a34.port_a_address_clear = "none";
defparam ram_block1a34.port_a_address_width = 13;
defparam ram_block1a34.port_a_byte_enable_mask_width = 1;
defparam ram_block1a34.port_a_byte_size = 1;
defparam ram_block1a34.port_a_data_out_clear = "none";
defparam ram_block1a34.port_a_data_out_clock = "none";
defparam ram_block1a34.port_a_data_width = 1;
defparam ram_block1a34.port_a_first_address = 0;
defparam ram_block1a34.port_a_first_bit_number = 34;
defparam ram_block1a34.port_a_last_address = 8191;
defparam ram_block1a34.port_a_logical_ram_depth = 16384;
defparam ram_block1a34.port_a_logical_ram_width = 64;
defparam ram_block1a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a34.port_b_address_clear = "none";
defparam ram_block1a34.port_b_address_clock = "clock1";
defparam ram_block1a34.port_b_address_width = 13;
defparam ram_block1a34.port_b_byte_enable_clock = "clock1";
defparam ram_block1a34.port_b_byte_enable_mask_width = 1;
defparam ram_block1a34.port_b_byte_size = 1;
defparam ram_block1a34.port_b_data_in_clock = "clock1";
defparam ram_block1a34.port_b_data_out_clear = "none";
defparam ram_block1a34.port_b_data_out_clock = "none";
defparam ram_block1a34.port_b_data_width = 1;
defparam ram_block1a34.port_b_first_address = 0;
defparam ram_block1a34.port_b_first_bit_number = 34;
defparam ram_block1a34.port_b_last_address = 8191;
defparam ram_block1a34.port_b_logical_ram_depth = 16384;
defparam ram_block1a34.port_b_logical_ram_width = 64;
defparam ram_block1a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a34.port_b_read_enable_clock = "clock1";
defparam ram_block1a34.port_b_write_enable_clock = "clock1";
defparam ram_block1a34.ram_block_type = "auto";
defparam ram_block1a34.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a34.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a34.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a34.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a99(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[35]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[35]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a99_PORTADATAOUT_bus),
	.portbdataout(ram_block1a99_PORTBDATAOUT_bus));
defparam ram_block1a99.clk0_core_clock_enable = "ena0";
defparam ram_block1a99.clk0_input_clock_enable = "ena0";
defparam ram_block1a99.clk1_core_clock_enable = "ena1";
defparam ram_block1a99.clk1_input_clock_enable = "ena1";
defparam ram_block1a99.data_interleave_offset_in_bits = 1;
defparam ram_block1a99.data_interleave_width_in_bits = 1;
defparam ram_block1a99.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a99.init_file_layout = "port_a";
defparam ram_block1a99.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a99.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a99.operation_mode = "bidir_dual_port";
defparam ram_block1a99.port_a_address_clear = "none";
defparam ram_block1a99.port_a_address_width = 13;
defparam ram_block1a99.port_a_byte_enable_mask_width = 1;
defparam ram_block1a99.port_a_byte_size = 1;
defparam ram_block1a99.port_a_data_out_clear = "none";
defparam ram_block1a99.port_a_data_out_clock = "none";
defparam ram_block1a99.port_a_data_width = 1;
defparam ram_block1a99.port_a_first_address = 8192;
defparam ram_block1a99.port_a_first_bit_number = 35;
defparam ram_block1a99.port_a_last_address = 16383;
defparam ram_block1a99.port_a_logical_ram_depth = 16384;
defparam ram_block1a99.port_a_logical_ram_width = 64;
defparam ram_block1a99.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a99.port_b_address_clear = "none";
defparam ram_block1a99.port_b_address_clock = "clock1";
defparam ram_block1a99.port_b_address_width = 13;
defparam ram_block1a99.port_b_byte_enable_clock = "clock1";
defparam ram_block1a99.port_b_byte_enable_mask_width = 1;
defparam ram_block1a99.port_b_byte_size = 1;
defparam ram_block1a99.port_b_data_in_clock = "clock1";
defparam ram_block1a99.port_b_data_out_clear = "none";
defparam ram_block1a99.port_b_data_out_clock = "none";
defparam ram_block1a99.port_b_data_width = 1;
defparam ram_block1a99.port_b_first_address = 8192;
defparam ram_block1a99.port_b_first_bit_number = 35;
defparam ram_block1a99.port_b_last_address = 16383;
defparam ram_block1a99.port_b_logical_ram_depth = 16384;
defparam ram_block1a99.port_b_logical_ram_width = 64;
defparam ram_block1a99.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a99.port_b_read_enable_clock = "clock1";
defparam ram_block1a99.port_b_write_enable_clock = "clock1";
defparam ram_block1a99.ram_block_type = "auto";
defparam ram_block1a99.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a99.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a99.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a99.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a35(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[35]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[35]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a35_PORTADATAOUT_bus),
	.portbdataout(ram_block1a35_PORTBDATAOUT_bus));
defparam ram_block1a35.clk0_core_clock_enable = "ena0";
defparam ram_block1a35.clk0_input_clock_enable = "ena0";
defparam ram_block1a35.clk1_core_clock_enable = "ena1";
defparam ram_block1a35.clk1_input_clock_enable = "ena1";
defparam ram_block1a35.data_interleave_offset_in_bits = 1;
defparam ram_block1a35.data_interleave_width_in_bits = 1;
defparam ram_block1a35.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a35.init_file_layout = "port_a";
defparam ram_block1a35.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a35.operation_mode = "bidir_dual_port";
defparam ram_block1a35.port_a_address_clear = "none";
defparam ram_block1a35.port_a_address_width = 13;
defparam ram_block1a35.port_a_byte_enable_mask_width = 1;
defparam ram_block1a35.port_a_byte_size = 1;
defparam ram_block1a35.port_a_data_out_clear = "none";
defparam ram_block1a35.port_a_data_out_clock = "none";
defparam ram_block1a35.port_a_data_width = 1;
defparam ram_block1a35.port_a_first_address = 0;
defparam ram_block1a35.port_a_first_bit_number = 35;
defparam ram_block1a35.port_a_last_address = 8191;
defparam ram_block1a35.port_a_logical_ram_depth = 16384;
defparam ram_block1a35.port_a_logical_ram_width = 64;
defparam ram_block1a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a35.port_b_address_clear = "none";
defparam ram_block1a35.port_b_address_clock = "clock1";
defparam ram_block1a35.port_b_address_width = 13;
defparam ram_block1a35.port_b_byte_enable_clock = "clock1";
defparam ram_block1a35.port_b_byte_enable_mask_width = 1;
defparam ram_block1a35.port_b_byte_size = 1;
defparam ram_block1a35.port_b_data_in_clock = "clock1";
defparam ram_block1a35.port_b_data_out_clear = "none";
defparam ram_block1a35.port_b_data_out_clock = "none";
defparam ram_block1a35.port_b_data_width = 1;
defparam ram_block1a35.port_b_first_address = 0;
defparam ram_block1a35.port_b_first_bit_number = 35;
defparam ram_block1a35.port_b_last_address = 8191;
defparam ram_block1a35.port_b_logical_ram_depth = 16384;
defparam ram_block1a35.port_b_logical_ram_width = 64;
defparam ram_block1a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a35.port_b_read_enable_clock = "clock1";
defparam ram_block1a35.port_b_write_enable_clock = "clock1";
defparam ram_block1a35.ram_block_type = "auto";
defparam ram_block1a35.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a35.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a35.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a35.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a100(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[36]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[36]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a100_PORTADATAOUT_bus),
	.portbdataout(ram_block1a100_PORTBDATAOUT_bus));
defparam ram_block1a100.clk0_core_clock_enable = "ena0";
defparam ram_block1a100.clk0_input_clock_enable = "ena0";
defparam ram_block1a100.clk1_core_clock_enable = "ena1";
defparam ram_block1a100.clk1_input_clock_enable = "ena1";
defparam ram_block1a100.data_interleave_offset_in_bits = 1;
defparam ram_block1a100.data_interleave_width_in_bits = 1;
defparam ram_block1a100.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a100.init_file_layout = "port_a";
defparam ram_block1a100.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a100.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a100.operation_mode = "bidir_dual_port";
defparam ram_block1a100.port_a_address_clear = "none";
defparam ram_block1a100.port_a_address_width = 13;
defparam ram_block1a100.port_a_byte_enable_mask_width = 1;
defparam ram_block1a100.port_a_byte_size = 1;
defparam ram_block1a100.port_a_data_out_clear = "none";
defparam ram_block1a100.port_a_data_out_clock = "none";
defparam ram_block1a100.port_a_data_width = 1;
defparam ram_block1a100.port_a_first_address = 8192;
defparam ram_block1a100.port_a_first_bit_number = 36;
defparam ram_block1a100.port_a_last_address = 16383;
defparam ram_block1a100.port_a_logical_ram_depth = 16384;
defparam ram_block1a100.port_a_logical_ram_width = 64;
defparam ram_block1a100.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a100.port_b_address_clear = "none";
defparam ram_block1a100.port_b_address_clock = "clock1";
defparam ram_block1a100.port_b_address_width = 13;
defparam ram_block1a100.port_b_byte_enable_clock = "clock1";
defparam ram_block1a100.port_b_byte_enable_mask_width = 1;
defparam ram_block1a100.port_b_byte_size = 1;
defparam ram_block1a100.port_b_data_in_clock = "clock1";
defparam ram_block1a100.port_b_data_out_clear = "none";
defparam ram_block1a100.port_b_data_out_clock = "none";
defparam ram_block1a100.port_b_data_width = 1;
defparam ram_block1a100.port_b_first_address = 8192;
defparam ram_block1a100.port_b_first_bit_number = 36;
defparam ram_block1a100.port_b_last_address = 16383;
defparam ram_block1a100.port_b_logical_ram_depth = 16384;
defparam ram_block1a100.port_b_logical_ram_width = 64;
defparam ram_block1a100.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a100.port_b_read_enable_clock = "clock1";
defparam ram_block1a100.port_b_write_enable_clock = "clock1";
defparam ram_block1a100.ram_block_type = "auto";
defparam ram_block1a100.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a100.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a100.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a100.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a36(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[36]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[36]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a36_PORTADATAOUT_bus),
	.portbdataout(ram_block1a36_PORTBDATAOUT_bus));
defparam ram_block1a36.clk0_core_clock_enable = "ena0";
defparam ram_block1a36.clk0_input_clock_enable = "ena0";
defparam ram_block1a36.clk1_core_clock_enable = "ena1";
defparam ram_block1a36.clk1_input_clock_enable = "ena1";
defparam ram_block1a36.data_interleave_offset_in_bits = 1;
defparam ram_block1a36.data_interleave_width_in_bits = 1;
defparam ram_block1a36.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a36.init_file_layout = "port_a";
defparam ram_block1a36.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a36.operation_mode = "bidir_dual_port";
defparam ram_block1a36.port_a_address_clear = "none";
defparam ram_block1a36.port_a_address_width = 13;
defparam ram_block1a36.port_a_byte_enable_mask_width = 1;
defparam ram_block1a36.port_a_byte_size = 1;
defparam ram_block1a36.port_a_data_out_clear = "none";
defparam ram_block1a36.port_a_data_out_clock = "none";
defparam ram_block1a36.port_a_data_width = 1;
defparam ram_block1a36.port_a_first_address = 0;
defparam ram_block1a36.port_a_first_bit_number = 36;
defparam ram_block1a36.port_a_last_address = 8191;
defparam ram_block1a36.port_a_logical_ram_depth = 16384;
defparam ram_block1a36.port_a_logical_ram_width = 64;
defparam ram_block1a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a36.port_b_address_clear = "none";
defparam ram_block1a36.port_b_address_clock = "clock1";
defparam ram_block1a36.port_b_address_width = 13;
defparam ram_block1a36.port_b_byte_enable_clock = "clock1";
defparam ram_block1a36.port_b_byte_enable_mask_width = 1;
defparam ram_block1a36.port_b_byte_size = 1;
defparam ram_block1a36.port_b_data_in_clock = "clock1";
defparam ram_block1a36.port_b_data_out_clear = "none";
defparam ram_block1a36.port_b_data_out_clock = "none";
defparam ram_block1a36.port_b_data_width = 1;
defparam ram_block1a36.port_b_first_address = 0;
defparam ram_block1a36.port_b_first_bit_number = 36;
defparam ram_block1a36.port_b_last_address = 8191;
defparam ram_block1a36.port_b_logical_ram_depth = 16384;
defparam ram_block1a36.port_b_logical_ram_width = 64;
defparam ram_block1a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a36.port_b_read_enable_clock = "clock1";
defparam ram_block1a36.port_b_write_enable_clock = "clock1";
defparam ram_block1a36.ram_block_type = "auto";
defparam ram_block1a36.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a36.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a36.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a36.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a101(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[37]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[37]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a101_PORTADATAOUT_bus),
	.portbdataout(ram_block1a101_PORTBDATAOUT_bus));
defparam ram_block1a101.clk0_core_clock_enable = "ena0";
defparam ram_block1a101.clk0_input_clock_enable = "ena0";
defparam ram_block1a101.clk1_core_clock_enable = "ena1";
defparam ram_block1a101.clk1_input_clock_enable = "ena1";
defparam ram_block1a101.data_interleave_offset_in_bits = 1;
defparam ram_block1a101.data_interleave_width_in_bits = 1;
defparam ram_block1a101.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a101.init_file_layout = "port_a";
defparam ram_block1a101.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a101.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a101.operation_mode = "bidir_dual_port";
defparam ram_block1a101.port_a_address_clear = "none";
defparam ram_block1a101.port_a_address_width = 13;
defparam ram_block1a101.port_a_byte_enable_mask_width = 1;
defparam ram_block1a101.port_a_byte_size = 1;
defparam ram_block1a101.port_a_data_out_clear = "none";
defparam ram_block1a101.port_a_data_out_clock = "none";
defparam ram_block1a101.port_a_data_width = 1;
defparam ram_block1a101.port_a_first_address = 8192;
defparam ram_block1a101.port_a_first_bit_number = 37;
defparam ram_block1a101.port_a_last_address = 16383;
defparam ram_block1a101.port_a_logical_ram_depth = 16384;
defparam ram_block1a101.port_a_logical_ram_width = 64;
defparam ram_block1a101.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a101.port_b_address_clear = "none";
defparam ram_block1a101.port_b_address_clock = "clock1";
defparam ram_block1a101.port_b_address_width = 13;
defparam ram_block1a101.port_b_byte_enable_clock = "clock1";
defparam ram_block1a101.port_b_byte_enable_mask_width = 1;
defparam ram_block1a101.port_b_byte_size = 1;
defparam ram_block1a101.port_b_data_in_clock = "clock1";
defparam ram_block1a101.port_b_data_out_clear = "none";
defparam ram_block1a101.port_b_data_out_clock = "none";
defparam ram_block1a101.port_b_data_width = 1;
defparam ram_block1a101.port_b_first_address = 8192;
defparam ram_block1a101.port_b_first_bit_number = 37;
defparam ram_block1a101.port_b_last_address = 16383;
defparam ram_block1a101.port_b_logical_ram_depth = 16384;
defparam ram_block1a101.port_b_logical_ram_width = 64;
defparam ram_block1a101.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a101.port_b_read_enable_clock = "clock1";
defparam ram_block1a101.port_b_write_enable_clock = "clock1";
defparam ram_block1a101.ram_block_type = "auto";
defparam ram_block1a101.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a101.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a101.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a101.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a37(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[37]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[37]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a37_PORTADATAOUT_bus),
	.portbdataout(ram_block1a37_PORTBDATAOUT_bus));
defparam ram_block1a37.clk0_core_clock_enable = "ena0";
defparam ram_block1a37.clk0_input_clock_enable = "ena0";
defparam ram_block1a37.clk1_core_clock_enable = "ena1";
defparam ram_block1a37.clk1_input_clock_enable = "ena1";
defparam ram_block1a37.data_interleave_offset_in_bits = 1;
defparam ram_block1a37.data_interleave_width_in_bits = 1;
defparam ram_block1a37.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a37.init_file_layout = "port_a";
defparam ram_block1a37.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a37.operation_mode = "bidir_dual_port";
defparam ram_block1a37.port_a_address_clear = "none";
defparam ram_block1a37.port_a_address_width = 13;
defparam ram_block1a37.port_a_byte_enable_mask_width = 1;
defparam ram_block1a37.port_a_byte_size = 1;
defparam ram_block1a37.port_a_data_out_clear = "none";
defparam ram_block1a37.port_a_data_out_clock = "none";
defparam ram_block1a37.port_a_data_width = 1;
defparam ram_block1a37.port_a_first_address = 0;
defparam ram_block1a37.port_a_first_bit_number = 37;
defparam ram_block1a37.port_a_last_address = 8191;
defparam ram_block1a37.port_a_logical_ram_depth = 16384;
defparam ram_block1a37.port_a_logical_ram_width = 64;
defparam ram_block1a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a37.port_b_address_clear = "none";
defparam ram_block1a37.port_b_address_clock = "clock1";
defparam ram_block1a37.port_b_address_width = 13;
defparam ram_block1a37.port_b_byte_enable_clock = "clock1";
defparam ram_block1a37.port_b_byte_enable_mask_width = 1;
defparam ram_block1a37.port_b_byte_size = 1;
defparam ram_block1a37.port_b_data_in_clock = "clock1";
defparam ram_block1a37.port_b_data_out_clear = "none";
defparam ram_block1a37.port_b_data_out_clock = "none";
defparam ram_block1a37.port_b_data_width = 1;
defparam ram_block1a37.port_b_first_address = 0;
defparam ram_block1a37.port_b_first_bit_number = 37;
defparam ram_block1a37.port_b_last_address = 8191;
defparam ram_block1a37.port_b_logical_ram_depth = 16384;
defparam ram_block1a37.port_b_logical_ram_width = 64;
defparam ram_block1a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a37.port_b_read_enable_clock = "clock1";
defparam ram_block1a37.port_b_write_enable_clock = "clock1";
defparam ram_block1a37.ram_block_type = "auto";
defparam ram_block1a37.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a37.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a37.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a37.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a102(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[38]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[38]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a102_PORTADATAOUT_bus),
	.portbdataout(ram_block1a102_PORTBDATAOUT_bus));
defparam ram_block1a102.clk0_core_clock_enable = "ena0";
defparam ram_block1a102.clk0_input_clock_enable = "ena0";
defparam ram_block1a102.clk1_core_clock_enable = "ena1";
defparam ram_block1a102.clk1_input_clock_enable = "ena1";
defparam ram_block1a102.data_interleave_offset_in_bits = 1;
defparam ram_block1a102.data_interleave_width_in_bits = 1;
defparam ram_block1a102.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a102.init_file_layout = "port_a";
defparam ram_block1a102.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a102.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a102.operation_mode = "bidir_dual_port";
defparam ram_block1a102.port_a_address_clear = "none";
defparam ram_block1a102.port_a_address_width = 13;
defparam ram_block1a102.port_a_byte_enable_mask_width = 1;
defparam ram_block1a102.port_a_byte_size = 1;
defparam ram_block1a102.port_a_data_out_clear = "none";
defparam ram_block1a102.port_a_data_out_clock = "none";
defparam ram_block1a102.port_a_data_width = 1;
defparam ram_block1a102.port_a_first_address = 8192;
defparam ram_block1a102.port_a_first_bit_number = 38;
defparam ram_block1a102.port_a_last_address = 16383;
defparam ram_block1a102.port_a_logical_ram_depth = 16384;
defparam ram_block1a102.port_a_logical_ram_width = 64;
defparam ram_block1a102.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a102.port_b_address_clear = "none";
defparam ram_block1a102.port_b_address_clock = "clock1";
defparam ram_block1a102.port_b_address_width = 13;
defparam ram_block1a102.port_b_byte_enable_clock = "clock1";
defparam ram_block1a102.port_b_byte_enable_mask_width = 1;
defparam ram_block1a102.port_b_byte_size = 1;
defparam ram_block1a102.port_b_data_in_clock = "clock1";
defparam ram_block1a102.port_b_data_out_clear = "none";
defparam ram_block1a102.port_b_data_out_clock = "none";
defparam ram_block1a102.port_b_data_width = 1;
defparam ram_block1a102.port_b_first_address = 8192;
defparam ram_block1a102.port_b_first_bit_number = 38;
defparam ram_block1a102.port_b_last_address = 16383;
defparam ram_block1a102.port_b_logical_ram_depth = 16384;
defparam ram_block1a102.port_b_logical_ram_width = 64;
defparam ram_block1a102.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a102.port_b_read_enable_clock = "clock1";
defparam ram_block1a102.port_b_write_enable_clock = "clock1";
defparam ram_block1a102.ram_block_type = "auto";
defparam ram_block1a102.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a102.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a102.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a102.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a38(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[38]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[38]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a38_PORTADATAOUT_bus),
	.portbdataout(ram_block1a38_PORTBDATAOUT_bus));
defparam ram_block1a38.clk0_core_clock_enable = "ena0";
defparam ram_block1a38.clk0_input_clock_enable = "ena0";
defparam ram_block1a38.clk1_core_clock_enable = "ena1";
defparam ram_block1a38.clk1_input_clock_enable = "ena1";
defparam ram_block1a38.data_interleave_offset_in_bits = 1;
defparam ram_block1a38.data_interleave_width_in_bits = 1;
defparam ram_block1a38.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a38.init_file_layout = "port_a";
defparam ram_block1a38.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a38.operation_mode = "bidir_dual_port";
defparam ram_block1a38.port_a_address_clear = "none";
defparam ram_block1a38.port_a_address_width = 13;
defparam ram_block1a38.port_a_byte_enable_mask_width = 1;
defparam ram_block1a38.port_a_byte_size = 1;
defparam ram_block1a38.port_a_data_out_clear = "none";
defparam ram_block1a38.port_a_data_out_clock = "none";
defparam ram_block1a38.port_a_data_width = 1;
defparam ram_block1a38.port_a_first_address = 0;
defparam ram_block1a38.port_a_first_bit_number = 38;
defparam ram_block1a38.port_a_last_address = 8191;
defparam ram_block1a38.port_a_logical_ram_depth = 16384;
defparam ram_block1a38.port_a_logical_ram_width = 64;
defparam ram_block1a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a38.port_b_address_clear = "none";
defparam ram_block1a38.port_b_address_clock = "clock1";
defparam ram_block1a38.port_b_address_width = 13;
defparam ram_block1a38.port_b_byte_enable_clock = "clock1";
defparam ram_block1a38.port_b_byte_enable_mask_width = 1;
defparam ram_block1a38.port_b_byte_size = 1;
defparam ram_block1a38.port_b_data_in_clock = "clock1";
defparam ram_block1a38.port_b_data_out_clear = "none";
defparam ram_block1a38.port_b_data_out_clock = "none";
defparam ram_block1a38.port_b_data_width = 1;
defparam ram_block1a38.port_b_first_address = 0;
defparam ram_block1a38.port_b_first_bit_number = 38;
defparam ram_block1a38.port_b_last_address = 8191;
defparam ram_block1a38.port_b_logical_ram_depth = 16384;
defparam ram_block1a38.port_b_logical_ram_width = 64;
defparam ram_block1a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a38.port_b_read_enable_clock = "clock1";
defparam ram_block1a38.port_b_write_enable_clock = "clock1";
defparam ram_block1a38.ram_block_type = "auto";
defparam ram_block1a38.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a38.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a38.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a38.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a103(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[39]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[39]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a103_PORTADATAOUT_bus),
	.portbdataout(ram_block1a103_PORTBDATAOUT_bus));
defparam ram_block1a103.clk0_core_clock_enable = "ena0";
defparam ram_block1a103.clk0_input_clock_enable = "ena0";
defparam ram_block1a103.clk1_core_clock_enable = "ena1";
defparam ram_block1a103.clk1_input_clock_enable = "ena1";
defparam ram_block1a103.data_interleave_offset_in_bits = 1;
defparam ram_block1a103.data_interleave_width_in_bits = 1;
defparam ram_block1a103.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a103.init_file_layout = "port_a";
defparam ram_block1a103.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a103.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a103.operation_mode = "bidir_dual_port";
defparam ram_block1a103.port_a_address_clear = "none";
defparam ram_block1a103.port_a_address_width = 13;
defparam ram_block1a103.port_a_byte_enable_mask_width = 1;
defparam ram_block1a103.port_a_byte_size = 1;
defparam ram_block1a103.port_a_data_out_clear = "none";
defparam ram_block1a103.port_a_data_out_clock = "none";
defparam ram_block1a103.port_a_data_width = 1;
defparam ram_block1a103.port_a_first_address = 8192;
defparam ram_block1a103.port_a_first_bit_number = 39;
defparam ram_block1a103.port_a_last_address = 16383;
defparam ram_block1a103.port_a_logical_ram_depth = 16384;
defparam ram_block1a103.port_a_logical_ram_width = 64;
defparam ram_block1a103.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a103.port_b_address_clear = "none";
defparam ram_block1a103.port_b_address_clock = "clock1";
defparam ram_block1a103.port_b_address_width = 13;
defparam ram_block1a103.port_b_byte_enable_clock = "clock1";
defparam ram_block1a103.port_b_byte_enable_mask_width = 1;
defparam ram_block1a103.port_b_byte_size = 1;
defparam ram_block1a103.port_b_data_in_clock = "clock1";
defparam ram_block1a103.port_b_data_out_clear = "none";
defparam ram_block1a103.port_b_data_out_clock = "none";
defparam ram_block1a103.port_b_data_width = 1;
defparam ram_block1a103.port_b_first_address = 8192;
defparam ram_block1a103.port_b_first_bit_number = 39;
defparam ram_block1a103.port_b_last_address = 16383;
defparam ram_block1a103.port_b_logical_ram_depth = 16384;
defparam ram_block1a103.port_b_logical_ram_width = 64;
defparam ram_block1a103.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a103.port_b_read_enable_clock = "clock1";
defparam ram_block1a103.port_b_write_enable_clock = "clock1";
defparam ram_block1a103.ram_block_type = "auto";
defparam ram_block1a103.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a103.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a103.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a103.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a39(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[39]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[4]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[39]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[4]}),
	.portadataout(ram_block1a39_PORTADATAOUT_bus),
	.portbdataout(ram_block1a39_PORTBDATAOUT_bus));
defparam ram_block1a39.clk0_core_clock_enable = "ena0";
defparam ram_block1a39.clk0_input_clock_enable = "ena0";
defparam ram_block1a39.clk1_core_clock_enable = "ena1";
defparam ram_block1a39.clk1_input_clock_enable = "ena1";
defparam ram_block1a39.data_interleave_offset_in_bits = 1;
defparam ram_block1a39.data_interleave_width_in_bits = 1;
defparam ram_block1a39.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a39.init_file_layout = "port_a";
defparam ram_block1a39.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a39.operation_mode = "bidir_dual_port";
defparam ram_block1a39.port_a_address_clear = "none";
defparam ram_block1a39.port_a_address_width = 13;
defparam ram_block1a39.port_a_byte_enable_mask_width = 1;
defparam ram_block1a39.port_a_byte_size = 1;
defparam ram_block1a39.port_a_data_out_clear = "none";
defparam ram_block1a39.port_a_data_out_clock = "none";
defparam ram_block1a39.port_a_data_width = 1;
defparam ram_block1a39.port_a_first_address = 0;
defparam ram_block1a39.port_a_first_bit_number = 39;
defparam ram_block1a39.port_a_last_address = 8191;
defparam ram_block1a39.port_a_logical_ram_depth = 16384;
defparam ram_block1a39.port_a_logical_ram_width = 64;
defparam ram_block1a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a39.port_b_address_clear = "none";
defparam ram_block1a39.port_b_address_clock = "clock1";
defparam ram_block1a39.port_b_address_width = 13;
defparam ram_block1a39.port_b_byte_enable_clock = "clock1";
defparam ram_block1a39.port_b_byte_enable_mask_width = 1;
defparam ram_block1a39.port_b_byte_size = 1;
defparam ram_block1a39.port_b_data_in_clock = "clock1";
defparam ram_block1a39.port_b_data_out_clear = "none";
defparam ram_block1a39.port_b_data_out_clock = "none";
defparam ram_block1a39.port_b_data_width = 1;
defparam ram_block1a39.port_b_first_address = 0;
defparam ram_block1a39.port_b_first_bit_number = 39;
defparam ram_block1a39.port_b_last_address = 8191;
defparam ram_block1a39.port_b_logical_ram_depth = 16384;
defparam ram_block1a39.port_b_logical_ram_width = 64;
defparam ram_block1a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a39.port_b_read_enable_clock = "clock1";
defparam ram_block1a39.port_b_write_enable_clock = "clock1";
defparam ram_block1a39.ram_block_type = "auto";
defparam ram_block1a39.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a39.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a39.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a39.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a104(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[40]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[40]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a104_PORTADATAOUT_bus),
	.portbdataout(ram_block1a104_PORTBDATAOUT_bus));
defparam ram_block1a104.clk0_core_clock_enable = "ena0";
defparam ram_block1a104.clk0_input_clock_enable = "ena0";
defparam ram_block1a104.clk1_core_clock_enable = "ena1";
defparam ram_block1a104.clk1_input_clock_enable = "ena1";
defparam ram_block1a104.data_interleave_offset_in_bits = 1;
defparam ram_block1a104.data_interleave_width_in_bits = 1;
defparam ram_block1a104.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a104.init_file_layout = "port_a";
defparam ram_block1a104.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a104.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a104.operation_mode = "bidir_dual_port";
defparam ram_block1a104.port_a_address_clear = "none";
defparam ram_block1a104.port_a_address_width = 13;
defparam ram_block1a104.port_a_byte_enable_mask_width = 1;
defparam ram_block1a104.port_a_byte_size = 1;
defparam ram_block1a104.port_a_data_out_clear = "none";
defparam ram_block1a104.port_a_data_out_clock = "none";
defparam ram_block1a104.port_a_data_width = 1;
defparam ram_block1a104.port_a_first_address = 8192;
defparam ram_block1a104.port_a_first_bit_number = 40;
defparam ram_block1a104.port_a_last_address = 16383;
defparam ram_block1a104.port_a_logical_ram_depth = 16384;
defparam ram_block1a104.port_a_logical_ram_width = 64;
defparam ram_block1a104.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a104.port_b_address_clear = "none";
defparam ram_block1a104.port_b_address_clock = "clock1";
defparam ram_block1a104.port_b_address_width = 13;
defparam ram_block1a104.port_b_byte_enable_clock = "clock1";
defparam ram_block1a104.port_b_byte_enable_mask_width = 1;
defparam ram_block1a104.port_b_byte_size = 1;
defparam ram_block1a104.port_b_data_in_clock = "clock1";
defparam ram_block1a104.port_b_data_out_clear = "none";
defparam ram_block1a104.port_b_data_out_clock = "none";
defparam ram_block1a104.port_b_data_width = 1;
defparam ram_block1a104.port_b_first_address = 8192;
defparam ram_block1a104.port_b_first_bit_number = 40;
defparam ram_block1a104.port_b_last_address = 16383;
defparam ram_block1a104.port_b_logical_ram_depth = 16384;
defparam ram_block1a104.port_b_logical_ram_width = 64;
defparam ram_block1a104.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a104.port_b_read_enable_clock = "clock1";
defparam ram_block1a104.port_b_write_enable_clock = "clock1";
defparam ram_block1a104.ram_block_type = "auto";
defparam ram_block1a104.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a104.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a104.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a104.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a40(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[40]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[40]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a40_PORTADATAOUT_bus),
	.portbdataout(ram_block1a40_PORTBDATAOUT_bus));
defparam ram_block1a40.clk0_core_clock_enable = "ena0";
defparam ram_block1a40.clk0_input_clock_enable = "ena0";
defparam ram_block1a40.clk1_core_clock_enable = "ena1";
defparam ram_block1a40.clk1_input_clock_enable = "ena1";
defparam ram_block1a40.data_interleave_offset_in_bits = 1;
defparam ram_block1a40.data_interleave_width_in_bits = 1;
defparam ram_block1a40.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a40.init_file_layout = "port_a";
defparam ram_block1a40.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a40.operation_mode = "bidir_dual_port";
defparam ram_block1a40.port_a_address_clear = "none";
defparam ram_block1a40.port_a_address_width = 13;
defparam ram_block1a40.port_a_byte_enable_mask_width = 1;
defparam ram_block1a40.port_a_byte_size = 1;
defparam ram_block1a40.port_a_data_out_clear = "none";
defparam ram_block1a40.port_a_data_out_clock = "none";
defparam ram_block1a40.port_a_data_width = 1;
defparam ram_block1a40.port_a_first_address = 0;
defparam ram_block1a40.port_a_first_bit_number = 40;
defparam ram_block1a40.port_a_last_address = 8191;
defparam ram_block1a40.port_a_logical_ram_depth = 16384;
defparam ram_block1a40.port_a_logical_ram_width = 64;
defparam ram_block1a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a40.port_b_address_clear = "none";
defparam ram_block1a40.port_b_address_clock = "clock1";
defparam ram_block1a40.port_b_address_width = 13;
defparam ram_block1a40.port_b_byte_enable_clock = "clock1";
defparam ram_block1a40.port_b_byte_enable_mask_width = 1;
defparam ram_block1a40.port_b_byte_size = 1;
defparam ram_block1a40.port_b_data_in_clock = "clock1";
defparam ram_block1a40.port_b_data_out_clear = "none";
defparam ram_block1a40.port_b_data_out_clock = "none";
defparam ram_block1a40.port_b_data_width = 1;
defparam ram_block1a40.port_b_first_address = 0;
defparam ram_block1a40.port_b_first_bit_number = 40;
defparam ram_block1a40.port_b_last_address = 8191;
defparam ram_block1a40.port_b_logical_ram_depth = 16384;
defparam ram_block1a40.port_b_logical_ram_width = 64;
defparam ram_block1a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a40.port_b_read_enable_clock = "clock1";
defparam ram_block1a40.port_b_write_enable_clock = "clock1";
defparam ram_block1a40.ram_block_type = "auto";
defparam ram_block1a40.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a40.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a40.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a40.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a105(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[41]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[41]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a105_PORTADATAOUT_bus),
	.portbdataout(ram_block1a105_PORTBDATAOUT_bus));
defparam ram_block1a105.clk0_core_clock_enable = "ena0";
defparam ram_block1a105.clk0_input_clock_enable = "ena0";
defparam ram_block1a105.clk1_core_clock_enable = "ena1";
defparam ram_block1a105.clk1_input_clock_enable = "ena1";
defparam ram_block1a105.data_interleave_offset_in_bits = 1;
defparam ram_block1a105.data_interleave_width_in_bits = 1;
defparam ram_block1a105.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a105.init_file_layout = "port_a";
defparam ram_block1a105.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a105.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a105.operation_mode = "bidir_dual_port";
defparam ram_block1a105.port_a_address_clear = "none";
defparam ram_block1a105.port_a_address_width = 13;
defparam ram_block1a105.port_a_byte_enable_mask_width = 1;
defparam ram_block1a105.port_a_byte_size = 1;
defparam ram_block1a105.port_a_data_out_clear = "none";
defparam ram_block1a105.port_a_data_out_clock = "none";
defparam ram_block1a105.port_a_data_width = 1;
defparam ram_block1a105.port_a_first_address = 8192;
defparam ram_block1a105.port_a_first_bit_number = 41;
defparam ram_block1a105.port_a_last_address = 16383;
defparam ram_block1a105.port_a_logical_ram_depth = 16384;
defparam ram_block1a105.port_a_logical_ram_width = 64;
defparam ram_block1a105.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a105.port_b_address_clear = "none";
defparam ram_block1a105.port_b_address_clock = "clock1";
defparam ram_block1a105.port_b_address_width = 13;
defparam ram_block1a105.port_b_byte_enable_clock = "clock1";
defparam ram_block1a105.port_b_byte_enable_mask_width = 1;
defparam ram_block1a105.port_b_byte_size = 1;
defparam ram_block1a105.port_b_data_in_clock = "clock1";
defparam ram_block1a105.port_b_data_out_clear = "none";
defparam ram_block1a105.port_b_data_out_clock = "none";
defparam ram_block1a105.port_b_data_width = 1;
defparam ram_block1a105.port_b_first_address = 8192;
defparam ram_block1a105.port_b_first_bit_number = 41;
defparam ram_block1a105.port_b_last_address = 16383;
defparam ram_block1a105.port_b_logical_ram_depth = 16384;
defparam ram_block1a105.port_b_logical_ram_width = 64;
defparam ram_block1a105.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a105.port_b_read_enable_clock = "clock1";
defparam ram_block1a105.port_b_write_enable_clock = "clock1";
defparam ram_block1a105.ram_block_type = "auto";
defparam ram_block1a105.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a105.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a105.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a105.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a41(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[41]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[41]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a41_PORTADATAOUT_bus),
	.portbdataout(ram_block1a41_PORTBDATAOUT_bus));
defparam ram_block1a41.clk0_core_clock_enable = "ena0";
defparam ram_block1a41.clk0_input_clock_enable = "ena0";
defparam ram_block1a41.clk1_core_clock_enable = "ena1";
defparam ram_block1a41.clk1_input_clock_enable = "ena1";
defparam ram_block1a41.data_interleave_offset_in_bits = 1;
defparam ram_block1a41.data_interleave_width_in_bits = 1;
defparam ram_block1a41.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a41.init_file_layout = "port_a";
defparam ram_block1a41.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a41.operation_mode = "bidir_dual_port";
defparam ram_block1a41.port_a_address_clear = "none";
defparam ram_block1a41.port_a_address_width = 13;
defparam ram_block1a41.port_a_byte_enable_mask_width = 1;
defparam ram_block1a41.port_a_byte_size = 1;
defparam ram_block1a41.port_a_data_out_clear = "none";
defparam ram_block1a41.port_a_data_out_clock = "none";
defparam ram_block1a41.port_a_data_width = 1;
defparam ram_block1a41.port_a_first_address = 0;
defparam ram_block1a41.port_a_first_bit_number = 41;
defparam ram_block1a41.port_a_last_address = 8191;
defparam ram_block1a41.port_a_logical_ram_depth = 16384;
defparam ram_block1a41.port_a_logical_ram_width = 64;
defparam ram_block1a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a41.port_b_address_clear = "none";
defparam ram_block1a41.port_b_address_clock = "clock1";
defparam ram_block1a41.port_b_address_width = 13;
defparam ram_block1a41.port_b_byte_enable_clock = "clock1";
defparam ram_block1a41.port_b_byte_enable_mask_width = 1;
defparam ram_block1a41.port_b_byte_size = 1;
defparam ram_block1a41.port_b_data_in_clock = "clock1";
defparam ram_block1a41.port_b_data_out_clear = "none";
defparam ram_block1a41.port_b_data_out_clock = "none";
defparam ram_block1a41.port_b_data_width = 1;
defparam ram_block1a41.port_b_first_address = 0;
defparam ram_block1a41.port_b_first_bit_number = 41;
defparam ram_block1a41.port_b_last_address = 8191;
defparam ram_block1a41.port_b_logical_ram_depth = 16384;
defparam ram_block1a41.port_b_logical_ram_width = 64;
defparam ram_block1a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a41.port_b_read_enable_clock = "clock1";
defparam ram_block1a41.port_b_write_enable_clock = "clock1";
defparam ram_block1a41.ram_block_type = "auto";
defparam ram_block1a41.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a41.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a41.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a41.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a106(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[42]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[42]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a106_PORTADATAOUT_bus),
	.portbdataout(ram_block1a106_PORTBDATAOUT_bus));
defparam ram_block1a106.clk0_core_clock_enable = "ena0";
defparam ram_block1a106.clk0_input_clock_enable = "ena0";
defparam ram_block1a106.clk1_core_clock_enable = "ena1";
defparam ram_block1a106.clk1_input_clock_enable = "ena1";
defparam ram_block1a106.data_interleave_offset_in_bits = 1;
defparam ram_block1a106.data_interleave_width_in_bits = 1;
defparam ram_block1a106.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a106.init_file_layout = "port_a";
defparam ram_block1a106.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a106.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a106.operation_mode = "bidir_dual_port";
defparam ram_block1a106.port_a_address_clear = "none";
defparam ram_block1a106.port_a_address_width = 13;
defparam ram_block1a106.port_a_byte_enable_mask_width = 1;
defparam ram_block1a106.port_a_byte_size = 1;
defparam ram_block1a106.port_a_data_out_clear = "none";
defparam ram_block1a106.port_a_data_out_clock = "none";
defparam ram_block1a106.port_a_data_width = 1;
defparam ram_block1a106.port_a_first_address = 8192;
defparam ram_block1a106.port_a_first_bit_number = 42;
defparam ram_block1a106.port_a_last_address = 16383;
defparam ram_block1a106.port_a_logical_ram_depth = 16384;
defparam ram_block1a106.port_a_logical_ram_width = 64;
defparam ram_block1a106.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a106.port_b_address_clear = "none";
defparam ram_block1a106.port_b_address_clock = "clock1";
defparam ram_block1a106.port_b_address_width = 13;
defparam ram_block1a106.port_b_byte_enable_clock = "clock1";
defparam ram_block1a106.port_b_byte_enable_mask_width = 1;
defparam ram_block1a106.port_b_byte_size = 1;
defparam ram_block1a106.port_b_data_in_clock = "clock1";
defparam ram_block1a106.port_b_data_out_clear = "none";
defparam ram_block1a106.port_b_data_out_clock = "none";
defparam ram_block1a106.port_b_data_width = 1;
defparam ram_block1a106.port_b_first_address = 8192;
defparam ram_block1a106.port_b_first_bit_number = 42;
defparam ram_block1a106.port_b_last_address = 16383;
defparam ram_block1a106.port_b_logical_ram_depth = 16384;
defparam ram_block1a106.port_b_logical_ram_width = 64;
defparam ram_block1a106.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a106.port_b_read_enable_clock = "clock1";
defparam ram_block1a106.port_b_write_enable_clock = "clock1";
defparam ram_block1a106.ram_block_type = "auto";
defparam ram_block1a106.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a106.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a106.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a106.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a42(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[42]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[42]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a42_PORTADATAOUT_bus),
	.portbdataout(ram_block1a42_PORTBDATAOUT_bus));
defparam ram_block1a42.clk0_core_clock_enable = "ena0";
defparam ram_block1a42.clk0_input_clock_enable = "ena0";
defparam ram_block1a42.clk1_core_clock_enable = "ena1";
defparam ram_block1a42.clk1_input_clock_enable = "ena1";
defparam ram_block1a42.data_interleave_offset_in_bits = 1;
defparam ram_block1a42.data_interleave_width_in_bits = 1;
defparam ram_block1a42.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a42.init_file_layout = "port_a";
defparam ram_block1a42.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a42.operation_mode = "bidir_dual_port";
defparam ram_block1a42.port_a_address_clear = "none";
defparam ram_block1a42.port_a_address_width = 13;
defparam ram_block1a42.port_a_byte_enable_mask_width = 1;
defparam ram_block1a42.port_a_byte_size = 1;
defparam ram_block1a42.port_a_data_out_clear = "none";
defparam ram_block1a42.port_a_data_out_clock = "none";
defparam ram_block1a42.port_a_data_width = 1;
defparam ram_block1a42.port_a_first_address = 0;
defparam ram_block1a42.port_a_first_bit_number = 42;
defparam ram_block1a42.port_a_last_address = 8191;
defparam ram_block1a42.port_a_logical_ram_depth = 16384;
defparam ram_block1a42.port_a_logical_ram_width = 64;
defparam ram_block1a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a42.port_b_address_clear = "none";
defparam ram_block1a42.port_b_address_clock = "clock1";
defparam ram_block1a42.port_b_address_width = 13;
defparam ram_block1a42.port_b_byte_enable_clock = "clock1";
defparam ram_block1a42.port_b_byte_enable_mask_width = 1;
defparam ram_block1a42.port_b_byte_size = 1;
defparam ram_block1a42.port_b_data_in_clock = "clock1";
defparam ram_block1a42.port_b_data_out_clear = "none";
defparam ram_block1a42.port_b_data_out_clock = "none";
defparam ram_block1a42.port_b_data_width = 1;
defparam ram_block1a42.port_b_first_address = 0;
defparam ram_block1a42.port_b_first_bit_number = 42;
defparam ram_block1a42.port_b_last_address = 8191;
defparam ram_block1a42.port_b_logical_ram_depth = 16384;
defparam ram_block1a42.port_b_logical_ram_width = 64;
defparam ram_block1a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a42.port_b_read_enable_clock = "clock1";
defparam ram_block1a42.port_b_write_enable_clock = "clock1";
defparam ram_block1a42.ram_block_type = "auto";
defparam ram_block1a42.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a42.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a42.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a42.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a107(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[43]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[43]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a107_PORTADATAOUT_bus),
	.portbdataout(ram_block1a107_PORTBDATAOUT_bus));
defparam ram_block1a107.clk0_core_clock_enable = "ena0";
defparam ram_block1a107.clk0_input_clock_enable = "ena0";
defparam ram_block1a107.clk1_core_clock_enable = "ena1";
defparam ram_block1a107.clk1_input_clock_enable = "ena1";
defparam ram_block1a107.data_interleave_offset_in_bits = 1;
defparam ram_block1a107.data_interleave_width_in_bits = 1;
defparam ram_block1a107.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a107.init_file_layout = "port_a";
defparam ram_block1a107.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a107.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a107.operation_mode = "bidir_dual_port";
defparam ram_block1a107.port_a_address_clear = "none";
defparam ram_block1a107.port_a_address_width = 13;
defparam ram_block1a107.port_a_byte_enable_mask_width = 1;
defparam ram_block1a107.port_a_byte_size = 1;
defparam ram_block1a107.port_a_data_out_clear = "none";
defparam ram_block1a107.port_a_data_out_clock = "none";
defparam ram_block1a107.port_a_data_width = 1;
defparam ram_block1a107.port_a_first_address = 8192;
defparam ram_block1a107.port_a_first_bit_number = 43;
defparam ram_block1a107.port_a_last_address = 16383;
defparam ram_block1a107.port_a_logical_ram_depth = 16384;
defparam ram_block1a107.port_a_logical_ram_width = 64;
defparam ram_block1a107.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a107.port_b_address_clear = "none";
defparam ram_block1a107.port_b_address_clock = "clock1";
defparam ram_block1a107.port_b_address_width = 13;
defparam ram_block1a107.port_b_byte_enable_clock = "clock1";
defparam ram_block1a107.port_b_byte_enable_mask_width = 1;
defparam ram_block1a107.port_b_byte_size = 1;
defparam ram_block1a107.port_b_data_in_clock = "clock1";
defparam ram_block1a107.port_b_data_out_clear = "none";
defparam ram_block1a107.port_b_data_out_clock = "none";
defparam ram_block1a107.port_b_data_width = 1;
defparam ram_block1a107.port_b_first_address = 8192;
defparam ram_block1a107.port_b_first_bit_number = 43;
defparam ram_block1a107.port_b_last_address = 16383;
defparam ram_block1a107.port_b_logical_ram_depth = 16384;
defparam ram_block1a107.port_b_logical_ram_width = 64;
defparam ram_block1a107.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a107.port_b_read_enable_clock = "clock1";
defparam ram_block1a107.port_b_write_enable_clock = "clock1";
defparam ram_block1a107.ram_block_type = "auto";
defparam ram_block1a107.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a107.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a107.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a107.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a43(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[43]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[43]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a43_PORTADATAOUT_bus),
	.portbdataout(ram_block1a43_PORTBDATAOUT_bus));
defparam ram_block1a43.clk0_core_clock_enable = "ena0";
defparam ram_block1a43.clk0_input_clock_enable = "ena0";
defparam ram_block1a43.clk1_core_clock_enable = "ena1";
defparam ram_block1a43.clk1_input_clock_enable = "ena1";
defparam ram_block1a43.data_interleave_offset_in_bits = 1;
defparam ram_block1a43.data_interleave_width_in_bits = 1;
defparam ram_block1a43.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a43.init_file_layout = "port_a";
defparam ram_block1a43.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a43.operation_mode = "bidir_dual_port";
defparam ram_block1a43.port_a_address_clear = "none";
defparam ram_block1a43.port_a_address_width = 13;
defparam ram_block1a43.port_a_byte_enable_mask_width = 1;
defparam ram_block1a43.port_a_byte_size = 1;
defparam ram_block1a43.port_a_data_out_clear = "none";
defparam ram_block1a43.port_a_data_out_clock = "none";
defparam ram_block1a43.port_a_data_width = 1;
defparam ram_block1a43.port_a_first_address = 0;
defparam ram_block1a43.port_a_first_bit_number = 43;
defparam ram_block1a43.port_a_last_address = 8191;
defparam ram_block1a43.port_a_logical_ram_depth = 16384;
defparam ram_block1a43.port_a_logical_ram_width = 64;
defparam ram_block1a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a43.port_b_address_clear = "none";
defparam ram_block1a43.port_b_address_clock = "clock1";
defparam ram_block1a43.port_b_address_width = 13;
defparam ram_block1a43.port_b_byte_enable_clock = "clock1";
defparam ram_block1a43.port_b_byte_enable_mask_width = 1;
defparam ram_block1a43.port_b_byte_size = 1;
defparam ram_block1a43.port_b_data_in_clock = "clock1";
defparam ram_block1a43.port_b_data_out_clear = "none";
defparam ram_block1a43.port_b_data_out_clock = "none";
defparam ram_block1a43.port_b_data_width = 1;
defparam ram_block1a43.port_b_first_address = 0;
defparam ram_block1a43.port_b_first_bit_number = 43;
defparam ram_block1a43.port_b_last_address = 8191;
defparam ram_block1a43.port_b_logical_ram_depth = 16384;
defparam ram_block1a43.port_b_logical_ram_width = 64;
defparam ram_block1a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a43.port_b_read_enable_clock = "clock1";
defparam ram_block1a43.port_b_write_enable_clock = "clock1";
defparam ram_block1a43.ram_block_type = "auto";
defparam ram_block1a43.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a43.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a43.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a43.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a108(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[44]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[44]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a108_PORTADATAOUT_bus),
	.portbdataout(ram_block1a108_PORTBDATAOUT_bus));
defparam ram_block1a108.clk0_core_clock_enable = "ena0";
defparam ram_block1a108.clk0_input_clock_enable = "ena0";
defparam ram_block1a108.clk1_core_clock_enable = "ena1";
defparam ram_block1a108.clk1_input_clock_enable = "ena1";
defparam ram_block1a108.data_interleave_offset_in_bits = 1;
defparam ram_block1a108.data_interleave_width_in_bits = 1;
defparam ram_block1a108.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a108.init_file_layout = "port_a";
defparam ram_block1a108.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a108.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a108.operation_mode = "bidir_dual_port";
defparam ram_block1a108.port_a_address_clear = "none";
defparam ram_block1a108.port_a_address_width = 13;
defparam ram_block1a108.port_a_byte_enable_mask_width = 1;
defparam ram_block1a108.port_a_byte_size = 1;
defparam ram_block1a108.port_a_data_out_clear = "none";
defparam ram_block1a108.port_a_data_out_clock = "none";
defparam ram_block1a108.port_a_data_width = 1;
defparam ram_block1a108.port_a_first_address = 8192;
defparam ram_block1a108.port_a_first_bit_number = 44;
defparam ram_block1a108.port_a_last_address = 16383;
defparam ram_block1a108.port_a_logical_ram_depth = 16384;
defparam ram_block1a108.port_a_logical_ram_width = 64;
defparam ram_block1a108.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a108.port_b_address_clear = "none";
defparam ram_block1a108.port_b_address_clock = "clock1";
defparam ram_block1a108.port_b_address_width = 13;
defparam ram_block1a108.port_b_byte_enable_clock = "clock1";
defparam ram_block1a108.port_b_byte_enable_mask_width = 1;
defparam ram_block1a108.port_b_byte_size = 1;
defparam ram_block1a108.port_b_data_in_clock = "clock1";
defparam ram_block1a108.port_b_data_out_clear = "none";
defparam ram_block1a108.port_b_data_out_clock = "none";
defparam ram_block1a108.port_b_data_width = 1;
defparam ram_block1a108.port_b_first_address = 8192;
defparam ram_block1a108.port_b_first_bit_number = 44;
defparam ram_block1a108.port_b_last_address = 16383;
defparam ram_block1a108.port_b_logical_ram_depth = 16384;
defparam ram_block1a108.port_b_logical_ram_width = 64;
defparam ram_block1a108.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a108.port_b_read_enable_clock = "clock1";
defparam ram_block1a108.port_b_write_enable_clock = "clock1";
defparam ram_block1a108.ram_block_type = "auto";
defparam ram_block1a108.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a108.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a108.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a108.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a44(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[44]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[44]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a44_PORTADATAOUT_bus),
	.portbdataout(ram_block1a44_PORTBDATAOUT_bus));
defparam ram_block1a44.clk0_core_clock_enable = "ena0";
defparam ram_block1a44.clk0_input_clock_enable = "ena0";
defparam ram_block1a44.clk1_core_clock_enable = "ena1";
defparam ram_block1a44.clk1_input_clock_enable = "ena1";
defparam ram_block1a44.data_interleave_offset_in_bits = 1;
defparam ram_block1a44.data_interleave_width_in_bits = 1;
defparam ram_block1a44.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a44.init_file_layout = "port_a";
defparam ram_block1a44.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a44.operation_mode = "bidir_dual_port";
defparam ram_block1a44.port_a_address_clear = "none";
defparam ram_block1a44.port_a_address_width = 13;
defparam ram_block1a44.port_a_byte_enable_mask_width = 1;
defparam ram_block1a44.port_a_byte_size = 1;
defparam ram_block1a44.port_a_data_out_clear = "none";
defparam ram_block1a44.port_a_data_out_clock = "none";
defparam ram_block1a44.port_a_data_width = 1;
defparam ram_block1a44.port_a_first_address = 0;
defparam ram_block1a44.port_a_first_bit_number = 44;
defparam ram_block1a44.port_a_last_address = 8191;
defparam ram_block1a44.port_a_logical_ram_depth = 16384;
defparam ram_block1a44.port_a_logical_ram_width = 64;
defparam ram_block1a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a44.port_b_address_clear = "none";
defparam ram_block1a44.port_b_address_clock = "clock1";
defparam ram_block1a44.port_b_address_width = 13;
defparam ram_block1a44.port_b_byte_enable_clock = "clock1";
defparam ram_block1a44.port_b_byte_enable_mask_width = 1;
defparam ram_block1a44.port_b_byte_size = 1;
defparam ram_block1a44.port_b_data_in_clock = "clock1";
defparam ram_block1a44.port_b_data_out_clear = "none";
defparam ram_block1a44.port_b_data_out_clock = "none";
defparam ram_block1a44.port_b_data_width = 1;
defparam ram_block1a44.port_b_first_address = 0;
defparam ram_block1a44.port_b_first_bit_number = 44;
defparam ram_block1a44.port_b_last_address = 8191;
defparam ram_block1a44.port_b_logical_ram_depth = 16384;
defparam ram_block1a44.port_b_logical_ram_width = 64;
defparam ram_block1a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a44.port_b_read_enable_clock = "clock1";
defparam ram_block1a44.port_b_write_enable_clock = "clock1";
defparam ram_block1a44.ram_block_type = "auto";
defparam ram_block1a44.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a44.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a44.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a44.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a109(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[45]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[45]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a109_PORTADATAOUT_bus),
	.portbdataout(ram_block1a109_PORTBDATAOUT_bus));
defparam ram_block1a109.clk0_core_clock_enable = "ena0";
defparam ram_block1a109.clk0_input_clock_enable = "ena0";
defparam ram_block1a109.clk1_core_clock_enable = "ena1";
defparam ram_block1a109.clk1_input_clock_enable = "ena1";
defparam ram_block1a109.data_interleave_offset_in_bits = 1;
defparam ram_block1a109.data_interleave_width_in_bits = 1;
defparam ram_block1a109.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a109.init_file_layout = "port_a";
defparam ram_block1a109.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a109.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a109.operation_mode = "bidir_dual_port";
defparam ram_block1a109.port_a_address_clear = "none";
defparam ram_block1a109.port_a_address_width = 13;
defparam ram_block1a109.port_a_byte_enable_mask_width = 1;
defparam ram_block1a109.port_a_byte_size = 1;
defparam ram_block1a109.port_a_data_out_clear = "none";
defparam ram_block1a109.port_a_data_out_clock = "none";
defparam ram_block1a109.port_a_data_width = 1;
defparam ram_block1a109.port_a_first_address = 8192;
defparam ram_block1a109.port_a_first_bit_number = 45;
defparam ram_block1a109.port_a_last_address = 16383;
defparam ram_block1a109.port_a_logical_ram_depth = 16384;
defparam ram_block1a109.port_a_logical_ram_width = 64;
defparam ram_block1a109.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a109.port_b_address_clear = "none";
defparam ram_block1a109.port_b_address_clock = "clock1";
defparam ram_block1a109.port_b_address_width = 13;
defparam ram_block1a109.port_b_byte_enable_clock = "clock1";
defparam ram_block1a109.port_b_byte_enable_mask_width = 1;
defparam ram_block1a109.port_b_byte_size = 1;
defparam ram_block1a109.port_b_data_in_clock = "clock1";
defparam ram_block1a109.port_b_data_out_clear = "none";
defparam ram_block1a109.port_b_data_out_clock = "none";
defparam ram_block1a109.port_b_data_width = 1;
defparam ram_block1a109.port_b_first_address = 8192;
defparam ram_block1a109.port_b_first_bit_number = 45;
defparam ram_block1a109.port_b_last_address = 16383;
defparam ram_block1a109.port_b_logical_ram_depth = 16384;
defparam ram_block1a109.port_b_logical_ram_width = 64;
defparam ram_block1a109.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a109.port_b_read_enable_clock = "clock1";
defparam ram_block1a109.port_b_write_enable_clock = "clock1";
defparam ram_block1a109.ram_block_type = "auto";
defparam ram_block1a109.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a109.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a109.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a109.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a45(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[45]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[45]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a45_PORTADATAOUT_bus),
	.portbdataout(ram_block1a45_PORTBDATAOUT_bus));
defparam ram_block1a45.clk0_core_clock_enable = "ena0";
defparam ram_block1a45.clk0_input_clock_enable = "ena0";
defparam ram_block1a45.clk1_core_clock_enable = "ena1";
defparam ram_block1a45.clk1_input_clock_enable = "ena1";
defparam ram_block1a45.data_interleave_offset_in_bits = 1;
defparam ram_block1a45.data_interleave_width_in_bits = 1;
defparam ram_block1a45.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a45.init_file_layout = "port_a";
defparam ram_block1a45.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a45.operation_mode = "bidir_dual_port";
defparam ram_block1a45.port_a_address_clear = "none";
defparam ram_block1a45.port_a_address_width = 13;
defparam ram_block1a45.port_a_byte_enable_mask_width = 1;
defparam ram_block1a45.port_a_byte_size = 1;
defparam ram_block1a45.port_a_data_out_clear = "none";
defparam ram_block1a45.port_a_data_out_clock = "none";
defparam ram_block1a45.port_a_data_width = 1;
defparam ram_block1a45.port_a_first_address = 0;
defparam ram_block1a45.port_a_first_bit_number = 45;
defparam ram_block1a45.port_a_last_address = 8191;
defparam ram_block1a45.port_a_logical_ram_depth = 16384;
defparam ram_block1a45.port_a_logical_ram_width = 64;
defparam ram_block1a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a45.port_b_address_clear = "none";
defparam ram_block1a45.port_b_address_clock = "clock1";
defparam ram_block1a45.port_b_address_width = 13;
defparam ram_block1a45.port_b_byte_enable_clock = "clock1";
defparam ram_block1a45.port_b_byte_enable_mask_width = 1;
defparam ram_block1a45.port_b_byte_size = 1;
defparam ram_block1a45.port_b_data_in_clock = "clock1";
defparam ram_block1a45.port_b_data_out_clear = "none";
defparam ram_block1a45.port_b_data_out_clock = "none";
defparam ram_block1a45.port_b_data_width = 1;
defparam ram_block1a45.port_b_first_address = 0;
defparam ram_block1a45.port_b_first_bit_number = 45;
defparam ram_block1a45.port_b_last_address = 8191;
defparam ram_block1a45.port_b_logical_ram_depth = 16384;
defparam ram_block1a45.port_b_logical_ram_width = 64;
defparam ram_block1a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a45.port_b_read_enable_clock = "clock1";
defparam ram_block1a45.port_b_write_enable_clock = "clock1";
defparam ram_block1a45.ram_block_type = "auto";
defparam ram_block1a45.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a45.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a45.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a45.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a110(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[46]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[46]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a110_PORTADATAOUT_bus),
	.portbdataout(ram_block1a110_PORTBDATAOUT_bus));
defparam ram_block1a110.clk0_core_clock_enable = "ena0";
defparam ram_block1a110.clk0_input_clock_enable = "ena0";
defparam ram_block1a110.clk1_core_clock_enable = "ena1";
defparam ram_block1a110.clk1_input_clock_enable = "ena1";
defparam ram_block1a110.data_interleave_offset_in_bits = 1;
defparam ram_block1a110.data_interleave_width_in_bits = 1;
defparam ram_block1a110.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a110.init_file_layout = "port_a";
defparam ram_block1a110.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a110.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a110.operation_mode = "bidir_dual_port";
defparam ram_block1a110.port_a_address_clear = "none";
defparam ram_block1a110.port_a_address_width = 13;
defparam ram_block1a110.port_a_byte_enable_mask_width = 1;
defparam ram_block1a110.port_a_byte_size = 1;
defparam ram_block1a110.port_a_data_out_clear = "none";
defparam ram_block1a110.port_a_data_out_clock = "none";
defparam ram_block1a110.port_a_data_width = 1;
defparam ram_block1a110.port_a_first_address = 8192;
defparam ram_block1a110.port_a_first_bit_number = 46;
defparam ram_block1a110.port_a_last_address = 16383;
defparam ram_block1a110.port_a_logical_ram_depth = 16384;
defparam ram_block1a110.port_a_logical_ram_width = 64;
defparam ram_block1a110.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a110.port_b_address_clear = "none";
defparam ram_block1a110.port_b_address_clock = "clock1";
defparam ram_block1a110.port_b_address_width = 13;
defparam ram_block1a110.port_b_byte_enable_clock = "clock1";
defparam ram_block1a110.port_b_byte_enable_mask_width = 1;
defparam ram_block1a110.port_b_byte_size = 1;
defparam ram_block1a110.port_b_data_in_clock = "clock1";
defparam ram_block1a110.port_b_data_out_clear = "none";
defparam ram_block1a110.port_b_data_out_clock = "none";
defparam ram_block1a110.port_b_data_width = 1;
defparam ram_block1a110.port_b_first_address = 8192;
defparam ram_block1a110.port_b_first_bit_number = 46;
defparam ram_block1a110.port_b_last_address = 16383;
defparam ram_block1a110.port_b_logical_ram_depth = 16384;
defparam ram_block1a110.port_b_logical_ram_width = 64;
defparam ram_block1a110.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a110.port_b_read_enable_clock = "clock1";
defparam ram_block1a110.port_b_write_enable_clock = "clock1";
defparam ram_block1a110.ram_block_type = "auto";
defparam ram_block1a110.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a110.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a110.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a110.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a46(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[46]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[46]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a46_PORTADATAOUT_bus),
	.portbdataout(ram_block1a46_PORTBDATAOUT_bus));
defparam ram_block1a46.clk0_core_clock_enable = "ena0";
defparam ram_block1a46.clk0_input_clock_enable = "ena0";
defparam ram_block1a46.clk1_core_clock_enable = "ena1";
defparam ram_block1a46.clk1_input_clock_enable = "ena1";
defparam ram_block1a46.data_interleave_offset_in_bits = 1;
defparam ram_block1a46.data_interleave_width_in_bits = 1;
defparam ram_block1a46.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a46.init_file_layout = "port_a";
defparam ram_block1a46.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a46.operation_mode = "bidir_dual_port";
defparam ram_block1a46.port_a_address_clear = "none";
defparam ram_block1a46.port_a_address_width = 13;
defparam ram_block1a46.port_a_byte_enable_mask_width = 1;
defparam ram_block1a46.port_a_byte_size = 1;
defparam ram_block1a46.port_a_data_out_clear = "none";
defparam ram_block1a46.port_a_data_out_clock = "none";
defparam ram_block1a46.port_a_data_width = 1;
defparam ram_block1a46.port_a_first_address = 0;
defparam ram_block1a46.port_a_first_bit_number = 46;
defparam ram_block1a46.port_a_last_address = 8191;
defparam ram_block1a46.port_a_logical_ram_depth = 16384;
defparam ram_block1a46.port_a_logical_ram_width = 64;
defparam ram_block1a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a46.port_b_address_clear = "none";
defparam ram_block1a46.port_b_address_clock = "clock1";
defparam ram_block1a46.port_b_address_width = 13;
defparam ram_block1a46.port_b_byte_enable_clock = "clock1";
defparam ram_block1a46.port_b_byte_enable_mask_width = 1;
defparam ram_block1a46.port_b_byte_size = 1;
defparam ram_block1a46.port_b_data_in_clock = "clock1";
defparam ram_block1a46.port_b_data_out_clear = "none";
defparam ram_block1a46.port_b_data_out_clock = "none";
defparam ram_block1a46.port_b_data_width = 1;
defparam ram_block1a46.port_b_first_address = 0;
defparam ram_block1a46.port_b_first_bit_number = 46;
defparam ram_block1a46.port_b_last_address = 8191;
defparam ram_block1a46.port_b_logical_ram_depth = 16384;
defparam ram_block1a46.port_b_logical_ram_width = 64;
defparam ram_block1a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a46.port_b_read_enable_clock = "clock1";
defparam ram_block1a46.port_b_write_enable_clock = "clock1";
defparam ram_block1a46.ram_block_type = "auto";
defparam ram_block1a46.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a46.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a46.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a46.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a111(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[47]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[47]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a111_PORTADATAOUT_bus),
	.portbdataout(ram_block1a111_PORTBDATAOUT_bus));
defparam ram_block1a111.clk0_core_clock_enable = "ena0";
defparam ram_block1a111.clk0_input_clock_enable = "ena0";
defparam ram_block1a111.clk1_core_clock_enable = "ena1";
defparam ram_block1a111.clk1_input_clock_enable = "ena1";
defparam ram_block1a111.data_interleave_offset_in_bits = 1;
defparam ram_block1a111.data_interleave_width_in_bits = 1;
defparam ram_block1a111.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a111.init_file_layout = "port_a";
defparam ram_block1a111.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a111.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a111.operation_mode = "bidir_dual_port";
defparam ram_block1a111.port_a_address_clear = "none";
defparam ram_block1a111.port_a_address_width = 13;
defparam ram_block1a111.port_a_byte_enable_mask_width = 1;
defparam ram_block1a111.port_a_byte_size = 1;
defparam ram_block1a111.port_a_data_out_clear = "none";
defparam ram_block1a111.port_a_data_out_clock = "none";
defparam ram_block1a111.port_a_data_width = 1;
defparam ram_block1a111.port_a_first_address = 8192;
defparam ram_block1a111.port_a_first_bit_number = 47;
defparam ram_block1a111.port_a_last_address = 16383;
defparam ram_block1a111.port_a_logical_ram_depth = 16384;
defparam ram_block1a111.port_a_logical_ram_width = 64;
defparam ram_block1a111.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a111.port_b_address_clear = "none";
defparam ram_block1a111.port_b_address_clock = "clock1";
defparam ram_block1a111.port_b_address_width = 13;
defparam ram_block1a111.port_b_byte_enable_clock = "clock1";
defparam ram_block1a111.port_b_byte_enable_mask_width = 1;
defparam ram_block1a111.port_b_byte_size = 1;
defparam ram_block1a111.port_b_data_in_clock = "clock1";
defparam ram_block1a111.port_b_data_out_clear = "none";
defparam ram_block1a111.port_b_data_out_clock = "none";
defparam ram_block1a111.port_b_data_width = 1;
defparam ram_block1a111.port_b_first_address = 8192;
defparam ram_block1a111.port_b_first_bit_number = 47;
defparam ram_block1a111.port_b_last_address = 16383;
defparam ram_block1a111.port_b_logical_ram_depth = 16384;
defparam ram_block1a111.port_b_logical_ram_width = 64;
defparam ram_block1a111.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a111.port_b_read_enable_clock = "clock1";
defparam ram_block1a111.port_b_write_enable_clock = "clock1";
defparam ram_block1a111.ram_block_type = "auto";
defparam ram_block1a111.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a111.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a111.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a111.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a47(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[47]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[5]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[47]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[5]}),
	.portadataout(ram_block1a47_PORTADATAOUT_bus),
	.portbdataout(ram_block1a47_PORTBDATAOUT_bus));
defparam ram_block1a47.clk0_core_clock_enable = "ena0";
defparam ram_block1a47.clk0_input_clock_enable = "ena0";
defparam ram_block1a47.clk1_core_clock_enable = "ena1";
defparam ram_block1a47.clk1_input_clock_enable = "ena1";
defparam ram_block1a47.data_interleave_offset_in_bits = 1;
defparam ram_block1a47.data_interleave_width_in_bits = 1;
defparam ram_block1a47.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a47.init_file_layout = "port_a";
defparam ram_block1a47.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a47.operation_mode = "bidir_dual_port";
defparam ram_block1a47.port_a_address_clear = "none";
defparam ram_block1a47.port_a_address_width = 13;
defparam ram_block1a47.port_a_byte_enable_mask_width = 1;
defparam ram_block1a47.port_a_byte_size = 1;
defparam ram_block1a47.port_a_data_out_clear = "none";
defparam ram_block1a47.port_a_data_out_clock = "none";
defparam ram_block1a47.port_a_data_width = 1;
defparam ram_block1a47.port_a_first_address = 0;
defparam ram_block1a47.port_a_first_bit_number = 47;
defparam ram_block1a47.port_a_last_address = 8191;
defparam ram_block1a47.port_a_logical_ram_depth = 16384;
defparam ram_block1a47.port_a_logical_ram_width = 64;
defparam ram_block1a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a47.port_b_address_clear = "none";
defparam ram_block1a47.port_b_address_clock = "clock1";
defparam ram_block1a47.port_b_address_width = 13;
defparam ram_block1a47.port_b_byte_enable_clock = "clock1";
defparam ram_block1a47.port_b_byte_enable_mask_width = 1;
defparam ram_block1a47.port_b_byte_size = 1;
defparam ram_block1a47.port_b_data_in_clock = "clock1";
defparam ram_block1a47.port_b_data_out_clear = "none";
defparam ram_block1a47.port_b_data_out_clock = "none";
defparam ram_block1a47.port_b_data_width = 1;
defparam ram_block1a47.port_b_first_address = 0;
defparam ram_block1a47.port_b_first_bit_number = 47;
defparam ram_block1a47.port_b_last_address = 8191;
defparam ram_block1a47.port_b_logical_ram_depth = 16384;
defparam ram_block1a47.port_b_logical_ram_width = 64;
defparam ram_block1a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a47.port_b_read_enable_clock = "clock1";
defparam ram_block1a47.port_b_write_enable_clock = "clock1";
defparam ram_block1a47.ram_block_type = "auto";
defparam ram_block1a47.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a47.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a47.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a47.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a112(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[48]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[48]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a112_PORTADATAOUT_bus),
	.portbdataout(ram_block1a112_PORTBDATAOUT_bus));
defparam ram_block1a112.clk0_core_clock_enable = "ena0";
defparam ram_block1a112.clk0_input_clock_enable = "ena0";
defparam ram_block1a112.clk1_core_clock_enable = "ena1";
defparam ram_block1a112.clk1_input_clock_enable = "ena1";
defparam ram_block1a112.data_interleave_offset_in_bits = 1;
defparam ram_block1a112.data_interleave_width_in_bits = 1;
defparam ram_block1a112.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a112.init_file_layout = "port_a";
defparam ram_block1a112.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a112.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a112.operation_mode = "bidir_dual_port";
defparam ram_block1a112.port_a_address_clear = "none";
defparam ram_block1a112.port_a_address_width = 13;
defparam ram_block1a112.port_a_byte_enable_mask_width = 1;
defparam ram_block1a112.port_a_byte_size = 1;
defparam ram_block1a112.port_a_data_out_clear = "none";
defparam ram_block1a112.port_a_data_out_clock = "none";
defparam ram_block1a112.port_a_data_width = 1;
defparam ram_block1a112.port_a_first_address = 8192;
defparam ram_block1a112.port_a_first_bit_number = 48;
defparam ram_block1a112.port_a_last_address = 16383;
defparam ram_block1a112.port_a_logical_ram_depth = 16384;
defparam ram_block1a112.port_a_logical_ram_width = 64;
defparam ram_block1a112.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a112.port_b_address_clear = "none";
defparam ram_block1a112.port_b_address_clock = "clock1";
defparam ram_block1a112.port_b_address_width = 13;
defparam ram_block1a112.port_b_byte_enable_clock = "clock1";
defparam ram_block1a112.port_b_byte_enable_mask_width = 1;
defparam ram_block1a112.port_b_byte_size = 1;
defparam ram_block1a112.port_b_data_in_clock = "clock1";
defparam ram_block1a112.port_b_data_out_clear = "none";
defparam ram_block1a112.port_b_data_out_clock = "none";
defparam ram_block1a112.port_b_data_width = 1;
defparam ram_block1a112.port_b_first_address = 8192;
defparam ram_block1a112.port_b_first_bit_number = 48;
defparam ram_block1a112.port_b_last_address = 16383;
defparam ram_block1a112.port_b_logical_ram_depth = 16384;
defparam ram_block1a112.port_b_logical_ram_width = 64;
defparam ram_block1a112.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a112.port_b_read_enable_clock = "clock1";
defparam ram_block1a112.port_b_write_enable_clock = "clock1";
defparam ram_block1a112.ram_block_type = "auto";
defparam ram_block1a112.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a112.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a112.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a112.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a48(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[48]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[48]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a48_PORTADATAOUT_bus),
	.portbdataout(ram_block1a48_PORTBDATAOUT_bus));
defparam ram_block1a48.clk0_core_clock_enable = "ena0";
defparam ram_block1a48.clk0_input_clock_enable = "ena0";
defparam ram_block1a48.clk1_core_clock_enable = "ena1";
defparam ram_block1a48.clk1_input_clock_enable = "ena1";
defparam ram_block1a48.data_interleave_offset_in_bits = 1;
defparam ram_block1a48.data_interleave_width_in_bits = 1;
defparam ram_block1a48.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a48.init_file_layout = "port_a";
defparam ram_block1a48.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a48.operation_mode = "bidir_dual_port";
defparam ram_block1a48.port_a_address_clear = "none";
defparam ram_block1a48.port_a_address_width = 13;
defparam ram_block1a48.port_a_byte_enable_mask_width = 1;
defparam ram_block1a48.port_a_byte_size = 1;
defparam ram_block1a48.port_a_data_out_clear = "none";
defparam ram_block1a48.port_a_data_out_clock = "none";
defparam ram_block1a48.port_a_data_width = 1;
defparam ram_block1a48.port_a_first_address = 0;
defparam ram_block1a48.port_a_first_bit_number = 48;
defparam ram_block1a48.port_a_last_address = 8191;
defparam ram_block1a48.port_a_logical_ram_depth = 16384;
defparam ram_block1a48.port_a_logical_ram_width = 64;
defparam ram_block1a48.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a48.port_b_address_clear = "none";
defparam ram_block1a48.port_b_address_clock = "clock1";
defparam ram_block1a48.port_b_address_width = 13;
defparam ram_block1a48.port_b_byte_enable_clock = "clock1";
defparam ram_block1a48.port_b_byte_enable_mask_width = 1;
defparam ram_block1a48.port_b_byte_size = 1;
defparam ram_block1a48.port_b_data_in_clock = "clock1";
defparam ram_block1a48.port_b_data_out_clear = "none";
defparam ram_block1a48.port_b_data_out_clock = "none";
defparam ram_block1a48.port_b_data_width = 1;
defparam ram_block1a48.port_b_first_address = 0;
defparam ram_block1a48.port_b_first_bit_number = 48;
defparam ram_block1a48.port_b_last_address = 8191;
defparam ram_block1a48.port_b_logical_ram_depth = 16384;
defparam ram_block1a48.port_b_logical_ram_width = 64;
defparam ram_block1a48.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a48.port_b_read_enable_clock = "clock1";
defparam ram_block1a48.port_b_write_enable_clock = "clock1";
defparam ram_block1a48.ram_block_type = "auto";
defparam ram_block1a48.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a48.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a48.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a48.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a113(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[49]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[49]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a113_PORTADATAOUT_bus),
	.portbdataout(ram_block1a113_PORTBDATAOUT_bus));
defparam ram_block1a113.clk0_core_clock_enable = "ena0";
defparam ram_block1a113.clk0_input_clock_enable = "ena0";
defparam ram_block1a113.clk1_core_clock_enable = "ena1";
defparam ram_block1a113.clk1_input_clock_enable = "ena1";
defparam ram_block1a113.data_interleave_offset_in_bits = 1;
defparam ram_block1a113.data_interleave_width_in_bits = 1;
defparam ram_block1a113.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a113.init_file_layout = "port_a";
defparam ram_block1a113.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a113.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a113.operation_mode = "bidir_dual_port";
defparam ram_block1a113.port_a_address_clear = "none";
defparam ram_block1a113.port_a_address_width = 13;
defparam ram_block1a113.port_a_byte_enable_mask_width = 1;
defparam ram_block1a113.port_a_byte_size = 1;
defparam ram_block1a113.port_a_data_out_clear = "none";
defparam ram_block1a113.port_a_data_out_clock = "none";
defparam ram_block1a113.port_a_data_width = 1;
defparam ram_block1a113.port_a_first_address = 8192;
defparam ram_block1a113.port_a_first_bit_number = 49;
defparam ram_block1a113.port_a_last_address = 16383;
defparam ram_block1a113.port_a_logical_ram_depth = 16384;
defparam ram_block1a113.port_a_logical_ram_width = 64;
defparam ram_block1a113.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a113.port_b_address_clear = "none";
defparam ram_block1a113.port_b_address_clock = "clock1";
defparam ram_block1a113.port_b_address_width = 13;
defparam ram_block1a113.port_b_byte_enable_clock = "clock1";
defparam ram_block1a113.port_b_byte_enable_mask_width = 1;
defparam ram_block1a113.port_b_byte_size = 1;
defparam ram_block1a113.port_b_data_in_clock = "clock1";
defparam ram_block1a113.port_b_data_out_clear = "none";
defparam ram_block1a113.port_b_data_out_clock = "none";
defparam ram_block1a113.port_b_data_width = 1;
defparam ram_block1a113.port_b_first_address = 8192;
defparam ram_block1a113.port_b_first_bit_number = 49;
defparam ram_block1a113.port_b_last_address = 16383;
defparam ram_block1a113.port_b_logical_ram_depth = 16384;
defparam ram_block1a113.port_b_logical_ram_width = 64;
defparam ram_block1a113.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a113.port_b_read_enable_clock = "clock1";
defparam ram_block1a113.port_b_write_enable_clock = "clock1";
defparam ram_block1a113.ram_block_type = "auto";
defparam ram_block1a113.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a113.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a113.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a113.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a49(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[49]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[49]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a49_PORTADATAOUT_bus),
	.portbdataout(ram_block1a49_PORTBDATAOUT_bus));
defparam ram_block1a49.clk0_core_clock_enable = "ena0";
defparam ram_block1a49.clk0_input_clock_enable = "ena0";
defparam ram_block1a49.clk1_core_clock_enable = "ena1";
defparam ram_block1a49.clk1_input_clock_enable = "ena1";
defparam ram_block1a49.data_interleave_offset_in_bits = 1;
defparam ram_block1a49.data_interleave_width_in_bits = 1;
defparam ram_block1a49.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a49.init_file_layout = "port_a";
defparam ram_block1a49.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a49.operation_mode = "bidir_dual_port";
defparam ram_block1a49.port_a_address_clear = "none";
defparam ram_block1a49.port_a_address_width = 13;
defparam ram_block1a49.port_a_byte_enable_mask_width = 1;
defparam ram_block1a49.port_a_byte_size = 1;
defparam ram_block1a49.port_a_data_out_clear = "none";
defparam ram_block1a49.port_a_data_out_clock = "none";
defparam ram_block1a49.port_a_data_width = 1;
defparam ram_block1a49.port_a_first_address = 0;
defparam ram_block1a49.port_a_first_bit_number = 49;
defparam ram_block1a49.port_a_last_address = 8191;
defparam ram_block1a49.port_a_logical_ram_depth = 16384;
defparam ram_block1a49.port_a_logical_ram_width = 64;
defparam ram_block1a49.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a49.port_b_address_clear = "none";
defparam ram_block1a49.port_b_address_clock = "clock1";
defparam ram_block1a49.port_b_address_width = 13;
defparam ram_block1a49.port_b_byte_enable_clock = "clock1";
defparam ram_block1a49.port_b_byte_enable_mask_width = 1;
defparam ram_block1a49.port_b_byte_size = 1;
defparam ram_block1a49.port_b_data_in_clock = "clock1";
defparam ram_block1a49.port_b_data_out_clear = "none";
defparam ram_block1a49.port_b_data_out_clock = "none";
defparam ram_block1a49.port_b_data_width = 1;
defparam ram_block1a49.port_b_first_address = 0;
defparam ram_block1a49.port_b_first_bit_number = 49;
defparam ram_block1a49.port_b_last_address = 8191;
defparam ram_block1a49.port_b_logical_ram_depth = 16384;
defparam ram_block1a49.port_b_logical_ram_width = 64;
defparam ram_block1a49.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a49.port_b_read_enable_clock = "clock1";
defparam ram_block1a49.port_b_write_enable_clock = "clock1";
defparam ram_block1a49.ram_block_type = "auto";
defparam ram_block1a49.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a49.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a49.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a49.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a114(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[50]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[50]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a114_PORTADATAOUT_bus),
	.portbdataout(ram_block1a114_PORTBDATAOUT_bus));
defparam ram_block1a114.clk0_core_clock_enable = "ena0";
defparam ram_block1a114.clk0_input_clock_enable = "ena0";
defparam ram_block1a114.clk1_core_clock_enable = "ena1";
defparam ram_block1a114.clk1_input_clock_enable = "ena1";
defparam ram_block1a114.data_interleave_offset_in_bits = 1;
defparam ram_block1a114.data_interleave_width_in_bits = 1;
defparam ram_block1a114.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a114.init_file_layout = "port_a";
defparam ram_block1a114.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a114.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a114.operation_mode = "bidir_dual_port";
defparam ram_block1a114.port_a_address_clear = "none";
defparam ram_block1a114.port_a_address_width = 13;
defparam ram_block1a114.port_a_byte_enable_mask_width = 1;
defparam ram_block1a114.port_a_byte_size = 1;
defparam ram_block1a114.port_a_data_out_clear = "none";
defparam ram_block1a114.port_a_data_out_clock = "none";
defparam ram_block1a114.port_a_data_width = 1;
defparam ram_block1a114.port_a_first_address = 8192;
defparam ram_block1a114.port_a_first_bit_number = 50;
defparam ram_block1a114.port_a_last_address = 16383;
defparam ram_block1a114.port_a_logical_ram_depth = 16384;
defparam ram_block1a114.port_a_logical_ram_width = 64;
defparam ram_block1a114.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a114.port_b_address_clear = "none";
defparam ram_block1a114.port_b_address_clock = "clock1";
defparam ram_block1a114.port_b_address_width = 13;
defparam ram_block1a114.port_b_byte_enable_clock = "clock1";
defparam ram_block1a114.port_b_byte_enable_mask_width = 1;
defparam ram_block1a114.port_b_byte_size = 1;
defparam ram_block1a114.port_b_data_in_clock = "clock1";
defparam ram_block1a114.port_b_data_out_clear = "none";
defparam ram_block1a114.port_b_data_out_clock = "none";
defparam ram_block1a114.port_b_data_width = 1;
defparam ram_block1a114.port_b_first_address = 8192;
defparam ram_block1a114.port_b_first_bit_number = 50;
defparam ram_block1a114.port_b_last_address = 16383;
defparam ram_block1a114.port_b_logical_ram_depth = 16384;
defparam ram_block1a114.port_b_logical_ram_width = 64;
defparam ram_block1a114.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a114.port_b_read_enable_clock = "clock1";
defparam ram_block1a114.port_b_write_enable_clock = "clock1";
defparam ram_block1a114.ram_block_type = "auto";
defparam ram_block1a114.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a114.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a114.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a114.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a50(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[50]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[50]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a50_PORTADATAOUT_bus),
	.portbdataout(ram_block1a50_PORTBDATAOUT_bus));
defparam ram_block1a50.clk0_core_clock_enable = "ena0";
defparam ram_block1a50.clk0_input_clock_enable = "ena0";
defparam ram_block1a50.clk1_core_clock_enable = "ena1";
defparam ram_block1a50.clk1_input_clock_enable = "ena1";
defparam ram_block1a50.data_interleave_offset_in_bits = 1;
defparam ram_block1a50.data_interleave_width_in_bits = 1;
defparam ram_block1a50.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a50.init_file_layout = "port_a";
defparam ram_block1a50.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a50.operation_mode = "bidir_dual_port";
defparam ram_block1a50.port_a_address_clear = "none";
defparam ram_block1a50.port_a_address_width = 13;
defparam ram_block1a50.port_a_byte_enable_mask_width = 1;
defparam ram_block1a50.port_a_byte_size = 1;
defparam ram_block1a50.port_a_data_out_clear = "none";
defparam ram_block1a50.port_a_data_out_clock = "none";
defparam ram_block1a50.port_a_data_width = 1;
defparam ram_block1a50.port_a_first_address = 0;
defparam ram_block1a50.port_a_first_bit_number = 50;
defparam ram_block1a50.port_a_last_address = 8191;
defparam ram_block1a50.port_a_logical_ram_depth = 16384;
defparam ram_block1a50.port_a_logical_ram_width = 64;
defparam ram_block1a50.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a50.port_b_address_clear = "none";
defparam ram_block1a50.port_b_address_clock = "clock1";
defparam ram_block1a50.port_b_address_width = 13;
defparam ram_block1a50.port_b_byte_enable_clock = "clock1";
defparam ram_block1a50.port_b_byte_enable_mask_width = 1;
defparam ram_block1a50.port_b_byte_size = 1;
defparam ram_block1a50.port_b_data_in_clock = "clock1";
defparam ram_block1a50.port_b_data_out_clear = "none";
defparam ram_block1a50.port_b_data_out_clock = "none";
defparam ram_block1a50.port_b_data_width = 1;
defparam ram_block1a50.port_b_first_address = 0;
defparam ram_block1a50.port_b_first_bit_number = 50;
defparam ram_block1a50.port_b_last_address = 8191;
defparam ram_block1a50.port_b_logical_ram_depth = 16384;
defparam ram_block1a50.port_b_logical_ram_width = 64;
defparam ram_block1a50.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a50.port_b_read_enable_clock = "clock1";
defparam ram_block1a50.port_b_write_enable_clock = "clock1";
defparam ram_block1a50.ram_block_type = "auto";
defparam ram_block1a50.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a50.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a50.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a50.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a115(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[51]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[51]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a115_PORTADATAOUT_bus),
	.portbdataout(ram_block1a115_PORTBDATAOUT_bus));
defparam ram_block1a115.clk0_core_clock_enable = "ena0";
defparam ram_block1a115.clk0_input_clock_enable = "ena0";
defparam ram_block1a115.clk1_core_clock_enable = "ena1";
defparam ram_block1a115.clk1_input_clock_enable = "ena1";
defparam ram_block1a115.data_interleave_offset_in_bits = 1;
defparam ram_block1a115.data_interleave_width_in_bits = 1;
defparam ram_block1a115.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a115.init_file_layout = "port_a";
defparam ram_block1a115.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a115.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a115.operation_mode = "bidir_dual_port";
defparam ram_block1a115.port_a_address_clear = "none";
defparam ram_block1a115.port_a_address_width = 13;
defparam ram_block1a115.port_a_byte_enable_mask_width = 1;
defparam ram_block1a115.port_a_byte_size = 1;
defparam ram_block1a115.port_a_data_out_clear = "none";
defparam ram_block1a115.port_a_data_out_clock = "none";
defparam ram_block1a115.port_a_data_width = 1;
defparam ram_block1a115.port_a_first_address = 8192;
defparam ram_block1a115.port_a_first_bit_number = 51;
defparam ram_block1a115.port_a_last_address = 16383;
defparam ram_block1a115.port_a_logical_ram_depth = 16384;
defparam ram_block1a115.port_a_logical_ram_width = 64;
defparam ram_block1a115.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a115.port_b_address_clear = "none";
defparam ram_block1a115.port_b_address_clock = "clock1";
defparam ram_block1a115.port_b_address_width = 13;
defparam ram_block1a115.port_b_byte_enable_clock = "clock1";
defparam ram_block1a115.port_b_byte_enable_mask_width = 1;
defparam ram_block1a115.port_b_byte_size = 1;
defparam ram_block1a115.port_b_data_in_clock = "clock1";
defparam ram_block1a115.port_b_data_out_clear = "none";
defparam ram_block1a115.port_b_data_out_clock = "none";
defparam ram_block1a115.port_b_data_width = 1;
defparam ram_block1a115.port_b_first_address = 8192;
defparam ram_block1a115.port_b_first_bit_number = 51;
defparam ram_block1a115.port_b_last_address = 16383;
defparam ram_block1a115.port_b_logical_ram_depth = 16384;
defparam ram_block1a115.port_b_logical_ram_width = 64;
defparam ram_block1a115.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a115.port_b_read_enable_clock = "clock1";
defparam ram_block1a115.port_b_write_enable_clock = "clock1";
defparam ram_block1a115.ram_block_type = "auto";
defparam ram_block1a115.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a115.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a115.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a115.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a51(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[51]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[51]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a51_PORTADATAOUT_bus),
	.portbdataout(ram_block1a51_PORTBDATAOUT_bus));
defparam ram_block1a51.clk0_core_clock_enable = "ena0";
defparam ram_block1a51.clk0_input_clock_enable = "ena0";
defparam ram_block1a51.clk1_core_clock_enable = "ena1";
defparam ram_block1a51.clk1_input_clock_enable = "ena1";
defparam ram_block1a51.data_interleave_offset_in_bits = 1;
defparam ram_block1a51.data_interleave_width_in_bits = 1;
defparam ram_block1a51.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a51.init_file_layout = "port_a";
defparam ram_block1a51.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a51.operation_mode = "bidir_dual_port";
defparam ram_block1a51.port_a_address_clear = "none";
defparam ram_block1a51.port_a_address_width = 13;
defparam ram_block1a51.port_a_byte_enable_mask_width = 1;
defparam ram_block1a51.port_a_byte_size = 1;
defparam ram_block1a51.port_a_data_out_clear = "none";
defparam ram_block1a51.port_a_data_out_clock = "none";
defparam ram_block1a51.port_a_data_width = 1;
defparam ram_block1a51.port_a_first_address = 0;
defparam ram_block1a51.port_a_first_bit_number = 51;
defparam ram_block1a51.port_a_last_address = 8191;
defparam ram_block1a51.port_a_logical_ram_depth = 16384;
defparam ram_block1a51.port_a_logical_ram_width = 64;
defparam ram_block1a51.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a51.port_b_address_clear = "none";
defparam ram_block1a51.port_b_address_clock = "clock1";
defparam ram_block1a51.port_b_address_width = 13;
defparam ram_block1a51.port_b_byte_enable_clock = "clock1";
defparam ram_block1a51.port_b_byte_enable_mask_width = 1;
defparam ram_block1a51.port_b_byte_size = 1;
defparam ram_block1a51.port_b_data_in_clock = "clock1";
defparam ram_block1a51.port_b_data_out_clear = "none";
defparam ram_block1a51.port_b_data_out_clock = "none";
defparam ram_block1a51.port_b_data_width = 1;
defparam ram_block1a51.port_b_first_address = 0;
defparam ram_block1a51.port_b_first_bit_number = 51;
defparam ram_block1a51.port_b_last_address = 8191;
defparam ram_block1a51.port_b_logical_ram_depth = 16384;
defparam ram_block1a51.port_b_logical_ram_width = 64;
defparam ram_block1a51.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a51.port_b_read_enable_clock = "clock1";
defparam ram_block1a51.port_b_write_enable_clock = "clock1";
defparam ram_block1a51.ram_block_type = "auto";
defparam ram_block1a51.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a51.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a51.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a51.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a116(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[52]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[52]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a116_PORTADATAOUT_bus),
	.portbdataout(ram_block1a116_PORTBDATAOUT_bus));
defparam ram_block1a116.clk0_core_clock_enable = "ena0";
defparam ram_block1a116.clk0_input_clock_enable = "ena0";
defparam ram_block1a116.clk1_core_clock_enable = "ena1";
defparam ram_block1a116.clk1_input_clock_enable = "ena1";
defparam ram_block1a116.data_interleave_offset_in_bits = 1;
defparam ram_block1a116.data_interleave_width_in_bits = 1;
defparam ram_block1a116.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a116.init_file_layout = "port_a";
defparam ram_block1a116.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a116.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a116.operation_mode = "bidir_dual_port";
defparam ram_block1a116.port_a_address_clear = "none";
defparam ram_block1a116.port_a_address_width = 13;
defparam ram_block1a116.port_a_byte_enable_mask_width = 1;
defparam ram_block1a116.port_a_byte_size = 1;
defparam ram_block1a116.port_a_data_out_clear = "none";
defparam ram_block1a116.port_a_data_out_clock = "none";
defparam ram_block1a116.port_a_data_width = 1;
defparam ram_block1a116.port_a_first_address = 8192;
defparam ram_block1a116.port_a_first_bit_number = 52;
defparam ram_block1a116.port_a_last_address = 16383;
defparam ram_block1a116.port_a_logical_ram_depth = 16384;
defparam ram_block1a116.port_a_logical_ram_width = 64;
defparam ram_block1a116.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a116.port_b_address_clear = "none";
defparam ram_block1a116.port_b_address_clock = "clock1";
defparam ram_block1a116.port_b_address_width = 13;
defparam ram_block1a116.port_b_byte_enable_clock = "clock1";
defparam ram_block1a116.port_b_byte_enable_mask_width = 1;
defparam ram_block1a116.port_b_byte_size = 1;
defparam ram_block1a116.port_b_data_in_clock = "clock1";
defparam ram_block1a116.port_b_data_out_clear = "none";
defparam ram_block1a116.port_b_data_out_clock = "none";
defparam ram_block1a116.port_b_data_width = 1;
defparam ram_block1a116.port_b_first_address = 8192;
defparam ram_block1a116.port_b_first_bit_number = 52;
defparam ram_block1a116.port_b_last_address = 16383;
defparam ram_block1a116.port_b_logical_ram_depth = 16384;
defparam ram_block1a116.port_b_logical_ram_width = 64;
defparam ram_block1a116.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a116.port_b_read_enable_clock = "clock1";
defparam ram_block1a116.port_b_write_enable_clock = "clock1";
defparam ram_block1a116.ram_block_type = "auto";
defparam ram_block1a116.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a116.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a116.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a116.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a52(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[52]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[52]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a52_PORTADATAOUT_bus),
	.portbdataout(ram_block1a52_PORTBDATAOUT_bus));
defparam ram_block1a52.clk0_core_clock_enable = "ena0";
defparam ram_block1a52.clk0_input_clock_enable = "ena0";
defparam ram_block1a52.clk1_core_clock_enable = "ena1";
defparam ram_block1a52.clk1_input_clock_enable = "ena1";
defparam ram_block1a52.data_interleave_offset_in_bits = 1;
defparam ram_block1a52.data_interleave_width_in_bits = 1;
defparam ram_block1a52.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a52.init_file_layout = "port_a";
defparam ram_block1a52.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a52.operation_mode = "bidir_dual_port";
defparam ram_block1a52.port_a_address_clear = "none";
defparam ram_block1a52.port_a_address_width = 13;
defparam ram_block1a52.port_a_byte_enable_mask_width = 1;
defparam ram_block1a52.port_a_byte_size = 1;
defparam ram_block1a52.port_a_data_out_clear = "none";
defparam ram_block1a52.port_a_data_out_clock = "none";
defparam ram_block1a52.port_a_data_width = 1;
defparam ram_block1a52.port_a_first_address = 0;
defparam ram_block1a52.port_a_first_bit_number = 52;
defparam ram_block1a52.port_a_last_address = 8191;
defparam ram_block1a52.port_a_logical_ram_depth = 16384;
defparam ram_block1a52.port_a_logical_ram_width = 64;
defparam ram_block1a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a52.port_b_address_clear = "none";
defparam ram_block1a52.port_b_address_clock = "clock1";
defparam ram_block1a52.port_b_address_width = 13;
defparam ram_block1a52.port_b_byte_enable_clock = "clock1";
defparam ram_block1a52.port_b_byte_enable_mask_width = 1;
defparam ram_block1a52.port_b_byte_size = 1;
defparam ram_block1a52.port_b_data_in_clock = "clock1";
defparam ram_block1a52.port_b_data_out_clear = "none";
defparam ram_block1a52.port_b_data_out_clock = "none";
defparam ram_block1a52.port_b_data_width = 1;
defparam ram_block1a52.port_b_first_address = 0;
defparam ram_block1a52.port_b_first_bit_number = 52;
defparam ram_block1a52.port_b_last_address = 8191;
defparam ram_block1a52.port_b_logical_ram_depth = 16384;
defparam ram_block1a52.port_b_logical_ram_width = 64;
defparam ram_block1a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a52.port_b_read_enable_clock = "clock1";
defparam ram_block1a52.port_b_write_enable_clock = "clock1";
defparam ram_block1a52.ram_block_type = "auto";
defparam ram_block1a52.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a52.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a52.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a52.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a117(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[53]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[53]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a117_PORTADATAOUT_bus),
	.portbdataout(ram_block1a117_PORTBDATAOUT_bus));
defparam ram_block1a117.clk0_core_clock_enable = "ena0";
defparam ram_block1a117.clk0_input_clock_enable = "ena0";
defparam ram_block1a117.clk1_core_clock_enable = "ena1";
defparam ram_block1a117.clk1_input_clock_enable = "ena1";
defparam ram_block1a117.data_interleave_offset_in_bits = 1;
defparam ram_block1a117.data_interleave_width_in_bits = 1;
defparam ram_block1a117.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a117.init_file_layout = "port_a";
defparam ram_block1a117.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a117.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a117.operation_mode = "bidir_dual_port";
defparam ram_block1a117.port_a_address_clear = "none";
defparam ram_block1a117.port_a_address_width = 13;
defparam ram_block1a117.port_a_byte_enable_mask_width = 1;
defparam ram_block1a117.port_a_byte_size = 1;
defparam ram_block1a117.port_a_data_out_clear = "none";
defparam ram_block1a117.port_a_data_out_clock = "none";
defparam ram_block1a117.port_a_data_width = 1;
defparam ram_block1a117.port_a_first_address = 8192;
defparam ram_block1a117.port_a_first_bit_number = 53;
defparam ram_block1a117.port_a_last_address = 16383;
defparam ram_block1a117.port_a_logical_ram_depth = 16384;
defparam ram_block1a117.port_a_logical_ram_width = 64;
defparam ram_block1a117.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a117.port_b_address_clear = "none";
defparam ram_block1a117.port_b_address_clock = "clock1";
defparam ram_block1a117.port_b_address_width = 13;
defparam ram_block1a117.port_b_byte_enable_clock = "clock1";
defparam ram_block1a117.port_b_byte_enable_mask_width = 1;
defparam ram_block1a117.port_b_byte_size = 1;
defparam ram_block1a117.port_b_data_in_clock = "clock1";
defparam ram_block1a117.port_b_data_out_clear = "none";
defparam ram_block1a117.port_b_data_out_clock = "none";
defparam ram_block1a117.port_b_data_width = 1;
defparam ram_block1a117.port_b_first_address = 8192;
defparam ram_block1a117.port_b_first_bit_number = 53;
defparam ram_block1a117.port_b_last_address = 16383;
defparam ram_block1a117.port_b_logical_ram_depth = 16384;
defparam ram_block1a117.port_b_logical_ram_width = 64;
defparam ram_block1a117.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a117.port_b_read_enable_clock = "clock1";
defparam ram_block1a117.port_b_write_enable_clock = "clock1";
defparam ram_block1a117.ram_block_type = "auto";
defparam ram_block1a117.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a117.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a117.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a117.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a53(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[53]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[53]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a53_PORTADATAOUT_bus),
	.portbdataout(ram_block1a53_PORTBDATAOUT_bus));
defparam ram_block1a53.clk0_core_clock_enable = "ena0";
defparam ram_block1a53.clk0_input_clock_enable = "ena0";
defparam ram_block1a53.clk1_core_clock_enable = "ena1";
defparam ram_block1a53.clk1_input_clock_enable = "ena1";
defparam ram_block1a53.data_interleave_offset_in_bits = 1;
defparam ram_block1a53.data_interleave_width_in_bits = 1;
defparam ram_block1a53.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a53.init_file_layout = "port_a";
defparam ram_block1a53.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a53.operation_mode = "bidir_dual_port";
defparam ram_block1a53.port_a_address_clear = "none";
defparam ram_block1a53.port_a_address_width = 13;
defparam ram_block1a53.port_a_byte_enable_mask_width = 1;
defparam ram_block1a53.port_a_byte_size = 1;
defparam ram_block1a53.port_a_data_out_clear = "none";
defparam ram_block1a53.port_a_data_out_clock = "none";
defparam ram_block1a53.port_a_data_width = 1;
defparam ram_block1a53.port_a_first_address = 0;
defparam ram_block1a53.port_a_first_bit_number = 53;
defparam ram_block1a53.port_a_last_address = 8191;
defparam ram_block1a53.port_a_logical_ram_depth = 16384;
defparam ram_block1a53.port_a_logical_ram_width = 64;
defparam ram_block1a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a53.port_b_address_clear = "none";
defparam ram_block1a53.port_b_address_clock = "clock1";
defparam ram_block1a53.port_b_address_width = 13;
defparam ram_block1a53.port_b_byte_enable_clock = "clock1";
defparam ram_block1a53.port_b_byte_enable_mask_width = 1;
defparam ram_block1a53.port_b_byte_size = 1;
defparam ram_block1a53.port_b_data_in_clock = "clock1";
defparam ram_block1a53.port_b_data_out_clear = "none";
defparam ram_block1a53.port_b_data_out_clock = "none";
defparam ram_block1a53.port_b_data_width = 1;
defparam ram_block1a53.port_b_first_address = 0;
defparam ram_block1a53.port_b_first_bit_number = 53;
defparam ram_block1a53.port_b_last_address = 8191;
defparam ram_block1a53.port_b_logical_ram_depth = 16384;
defparam ram_block1a53.port_b_logical_ram_width = 64;
defparam ram_block1a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a53.port_b_read_enable_clock = "clock1";
defparam ram_block1a53.port_b_write_enable_clock = "clock1";
defparam ram_block1a53.ram_block_type = "auto";
defparam ram_block1a53.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a53.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a53.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a53.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a118(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[54]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[54]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a118_PORTADATAOUT_bus),
	.portbdataout(ram_block1a118_PORTBDATAOUT_bus));
defparam ram_block1a118.clk0_core_clock_enable = "ena0";
defparam ram_block1a118.clk0_input_clock_enable = "ena0";
defparam ram_block1a118.clk1_core_clock_enable = "ena1";
defparam ram_block1a118.clk1_input_clock_enable = "ena1";
defparam ram_block1a118.data_interleave_offset_in_bits = 1;
defparam ram_block1a118.data_interleave_width_in_bits = 1;
defparam ram_block1a118.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a118.init_file_layout = "port_a";
defparam ram_block1a118.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a118.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a118.operation_mode = "bidir_dual_port";
defparam ram_block1a118.port_a_address_clear = "none";
defparam ram_block1a118.port_a_address_width = 13;
defparam ram_block1a118.port_a_byte_enable_mask_width = 1;
defparam ram_block1a118.port_a_byte_size = 1;
defparam ram_block1a118.port_a_data_out_clear = "none";
defparam ram_block1a118.port_a_data_out_clock = "none";
defparam ram_block1a118.port_a_data_width = 1;
defparam ram_block1a118.port_a_first_address = 8192;
defparam ram_block1a118.port_a_first_bit_number = 54;
defparam ram_block1a118.port_a_last_address = 16383;
defparam ram_block1a118.port_a_logical_ram_depth = 16384;
defparam ram_block1a118.port_a_logical_ram_width = 64;
defparam ram_block1a118.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a118.port_b_address_clear = "none";
defparam ram_block1a118.port_b_address_clock = "clock1";
defparam ram_block1a118.port_b_address_width = 13;
defparam ram_block1a118.port_b_byte_enable_clock = "clock1";
defparam ram_block1a118.port_b_byte_enable_mask_width = 1;
defparam ram_block1a118.port_b_byte_size = 1;
defparam ram_block1a118.port_b_data_in_clock = "clock1";
defparam ram_block1a118.port_b_data_out_clear = "none";
defparam ram_block1a118.port_b_data_out_clock = "none";
defparam ram_block1a118.port_b_data_width = 1;
defparam ram_block1a118.port_b_first_address = 8192;
defparam ram_block1a118.port_b_first_bit_number = 54;
defparam ram_block1a118.port_b_last_address = 16383;
defparam ram_block1a118.port_b_logical_ram_depth = 16384;
defparam ram_block1a118.port_b_logical_ram_width = 64;
defparam ram_block1a118.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a118.port_b_read_enable_clock = "clock1";
defparam ram_block1a118.port_b_write_enable_clock = "clock1";
defparam ram_block1a118.ram_block_type = "auto";
defparam ram_block1a118.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a118.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a118.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a118.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a54(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[54]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[54]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a54_PORTADATAOUT_bus),
	.portbdataout(ram_block1a54_PORTBDATAOUT_bus));
defparam ram_block1a54.clk0_core_clock_enable = "ena0";
defparam ram_block1a54.clk0_input_clock_enable = "ena0";
defparam ram_block1a54.clk1_core_clock_enable = "ena1";
defparam ram_block1a54.clk1_input_clock_enable = "ena1";
defparam ram_block1a54.data_interleave_offset_in_bits = 1;
defparam ram_block1a54.data_interleave_width_in_bits = 1;
defparam ram_block1a54.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a54.init_file_layout = "port_a";
defparam ram_block1a54.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a54.operation_mode = "bidir_dual_port";
defparam ram_block1a54.port_a_address_clear = "none";
defparam ram_block1a54.port_a_address_width = 13;
defparam ram_block1a54.port_a_byte_enable_mask_width = 1;
defparam ram_block1a54.port_a_byte_size = 1;
defparam ram_block1a54.port_a_data_out_clear = "none";
defparam ram_block1a54.port_a_data_out_clock = "none";
defparam ram_block1a54.port_a_data_width = 1;
defparam ram_block1a54.port_a_first_address = 0;
defparam ram_block1a54.port_a_first_bit_number = 54;
defparam ram_block1a54.port_a_last_address = 8191;
defparam ram_block1a54.port_a_logical_ram_depth = 16384;
defparam ram_block1a54.port_a_logical_ram_width = 64;
defparam ram_block1a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a54.port_b_address_clear = "none";
defparam ram_block1a54.port_b_address_clock = "clock1";
defparam ram_block1a54.port_b_address_width = 13;
defparam ram_block1a54.port_b_byte_enable_clock = "clock1";
defparam ram_block1a54.port_b_byte_enable_mask_width = 1;
defparam ram_block1a54.port_b_byte_size = 1;
defparam ram_block1a54.port_b_data_in_clock = "clock1";
defparam ram_block1a54.port_b_data_out_clear = "none";
defparam ram_block1a54.port_b_data_out_clock = "none";
defparam ram_block1a54.port_b_data_width = 1;
defparam ram_block1a54.port_b_first_address = 0;
defparam ram_block1a54.port_b_first_bit_number = 54;
defparam ram_block1a54.port_b_last_address = 8191;
defparam ram_block1a54.port_b_logical_ram_depth = 16384;
defparam ram_block1a54.port_b_logical_ram_width = 64;
defparam ram_block1a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a54.port_b_read_enable_clock = "clock1";
defparam ram_block1a54.port_b_write_enable_clock = "clock1";
defparam ram_block1a54.ram_block_type = "auto";
defparam ram_block1a54.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a54.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a54.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a54.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a119(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[55]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[55]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a119_PORTADATAOUT_bus),
	.portbdataout(ram_block1a119_PORTBDATAOUT_bus));
defparam ram_block1a119.clk0_core_clock_enable = "ena0";
defparam ram_block1a119.clk0_input_clock_enable = "ena0";
defparam ram_block1a119.clk1_core_clock_enable = "ena1";
defparam ram_block1a119.clk1_input_clock_enable = "ena1";
defparam ram_block1a119.data_interleave_offset_in_bits = 1;
defparam ram_block1a119.data_interleave_width_in_bits = 1;
defparam ram_block1a119.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a119.init_file_layout = "port_a";
defparam ram_block1a119.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a119.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a119.operation_mode = "bidir_dual_port";
defparam ram_block1a119.port_a_address_clear = "none";
defparam ram_block1a119.port_a_address_width = 13;
defparam ram_block1a119.port_a_byte_enable_mask_width = 1;
defparam ram_block1a119.port_a_byte_size = 1;
defparam ram_block1a119.port_a_data_out_clear = "none";
defparam ram_block1a119.port_a_data_out_clock = "none";
defparam ram_block1a119.port_a_data_width = 1;
defparam ram_block1a119.port_a_first_address = 8192;
defparam ram_block1a119.port_a_first_bit_number = 55;
defparam ram_block1a119.port_a_last_address = 16383;
defparam ram_block1a119.port_a_logical_ram_depth = 16384;
defparam ram_block1a119.port_a_logical_ram_width = 64;
defparam ram_block1a119.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a119.port_b_address_clear = "none";
defparam ram_block1a119.port_b_address_clock = "clock1";
defparam ram_block1a119.port_b_address_width = 13;
defparam ram_block1a119.port_b_byte_enable_clock = "clock1";
defparam ram_block1a119.port_b_byte_enable_mask_width = 1;
defparam ram_block1a119.port_b_byte_size = 1;
defparam ram_block1a119.port_b_data_in_clock = "clock1";
defparam ram_block1a119.port_b_data_out_clear = "none";
defparam ram_block1a119.port_b_data_out_clock = "none";
defparam ram_block1a119.port_b_data_width = 1;
defparam ram_block1a119.port_b_first_address = 8192;
defparam ram_block1a119.port_b_first_bit_number = 55;
defparam ram_block1a119.port_b_last_address = 16383;
defparam ram_block1a119.port_b_logical_ram_depth = 16384;
defparam ram_block1a119.port_b_logical_ram_width = 64;
defparam ram_block1a119.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a119.port_b_read_enable_clock = "clock1";
defparam ram_block1a119.port_b_write_enable_clock = "clock1";
defparam ram_block1a119.ram_block_type = "auto";
defparam ram_block1a119.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a119.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a119.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a119.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a55(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[55]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[6]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[55]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[6]}),
	.portadataout(ram_block1a55_PORTADATAOUT_bus),
	.portbdataout(ram_block1a55_PORTBDATAOUT_bus));
defparam ram_block1a55.clk0_core_clock_enable = "ena0";
defparam ram_block1a55.clk0_input_clock_enable = "ena0";
defparam ram_block1a55.clk1_core_clock_enable = "ena1";
defparam ram_block1a55.clk1_input_clock_enable = "ena1";
defparam ram_block1a55.data_interleave_offset_in_bits = 1;
defparam ram_block1a55.data_interleave_width_in_bits = 1;
defparam ram_block1a55.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a55.init_file_layout = "port_a";
defparam ram_block1a55.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a55.operation_mode = "bidir_dual_port";
defparam ram_block1a55.port_a_address_clear = "none";
defparam ram_block1a55.port_a_address_width = 13;
defparam ram_block1a55.port_a_byte_enable_mask_width = 1;
defparam ram_block1a55.port_a_byte_size = 1;
defparam ram_block1a55.port_a_data_out_clear = "none";
defparam ram_block1a55.port_a_data_out_clock = "none";
defparam ram_block1a55.port_a_data_width = 1;
defparam ram_block1a55.port_a_first_address = 0;
defparam ram_block1a55.port_a_first_bit_number = 55;
defparam ram_block1a55.port_a_last_address = 8191;
defparam ram_block1a55.port_a_logical_ram_depth = 16384;
defparam ram_block1a55.port_a_logical_ram_width = 64;
defparam ram_block1a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a55.port_b_address_clear = "none";
defparam ram_block1a55.port_b_address_clock = "clock1";
defparam ram_block1a55.port_b_address_width = 13;
defparam ram_block1a55.port_b_byte_enable_clock = "clock1";
defparam ram_block1a55.port_b_byte_enable_mask_width = 1;
defparam ram_block1a55.port_b_byte_size = 1;
defparam ram_block1a55.port_b_data_in_clock = "clock1";
defparam ram_block1a55.port_b_data_out_clear = "none";
defparam ram_block1a55.port_b_data_out_clock = "none";
defparam ram_block1a55.port_b_data_width = 1;
defparam ram_block1a55.port_b_first_address = 0;
defparam ram_block1a55.port_b_first_bit_number = 55;
defparam ram_block1a55.port_b_last_address = 8191;
defparam ram_block1a55.port_b_logical_ram_depth = 16384;
defparam ram_block1a55.port_b_logical_ram_width = 64;
defparam ram_block1a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a55.port_b_read_enable_clock = "clock1";
defparam ram_block1a55.port_b_write_enable_clock = "clock1";
defparam ram_block1a55.ram_block_type = "auto";
defparam ram_block1a55.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a55.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a55.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a55.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a120(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[56]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[56]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a120_PORTADATAOUT_bus),
	.portbdataout(ram_block1a120_PORTBDATAOUT_bus));
defparam ram_block1a120.clk0_core_clock_enable = "ena0";
defparam ram_block1a120.clk0_input_clock_enable = "ena0";
defparam ram_block1a120.clk1_core_clock_enable = "ena1";
defparam ram_block1a120.clk1_input_clock_enable = "ena1";
defparam ram_block1a120.data_interleave_offset_in_bits = 1;
defparam ram_block1a120.data_interleave_width_in_bits = 1;
defparam ram_block1a120.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a120.init_file_layout = "port_a";
defparam ram_block1a120.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a120.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a120.operation_mode = "bidir_dual_port";
defparam ram_block1a120.port_a_address_clear = "none";
defparam ram_block1a120.port_a_address_width = 13;
defparam ram_block1a120.port_a_byte_enable_mask_width = 1;
defparam ram_block1a120.port_a_byte_size = 1;
defparam ram_block1a120.port_a_data_out_clear = "none";
defparam ram_block1a120.port_a_data_out_clock = "none";
defparam ram_block1a120.port_a_data_width = 1;
defparam ram_block1a120.port_a_first_address = 8192;
defparam ram_block1a120.port_a_first_bit_number = 56;
defparam ram_block1a120.port_a_last_address = 16383;
defparam ram_block1a120.port_a_logical_ram_depth = 16384;
defparam ram_block1a120.port_a_logical_ram_width = 64;
defparam ram_block1a120.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a120.port_b_address_clear = "none";
defparam ram_block1a120.port_b_address_clock = "clock1";
defparam ram_block1a120.port_b_address_width = 13;
defparam ram_block1a120.port_b_byte_enable_clock = "clock1";
defparam ram_block1a120.port_b_byte_enable_mask_width = 1;
defparam ram_block1a120.port_b_byte_size = 1;
defparam ram_block1a120.port_b_data_in_clock = "clock1";
defparam ram_block1a120.port_b_data_out_clear = "none";
defparam ram_block1a120.port_b_data_out_clock = "none";
defparam ram_block1a120.port_b_data_width = 1;
defparam ram_block1a120.port_b_first_address = 8192;
defparam ram_block1a120.port_b_first_bit_number = 56;
defparam ram_block1a120.port_b_last_address = 16383;
defparam ram_block1a120.port_b_logical_ram_depth = 16384;
defparam ram_block1a120.port_b_logical_ram_width = 64;
defparam ram_block1a120.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a120.port_b_read_enable_clock = "clock1";
defparam ram_block1a120.port_b_write_enable_clock = "clock1";
defparam ram_block1a120.ram_block_type = "auto";
defparam ram_block1a120.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a120.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a120.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a120.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a56(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[56]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[56]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a56_PORTADATAOUT_bus),
	.portbdataout(ram_block1a56_PORTBDATAOUT_bus));
defparam ram_block1a56.clk0_core_clock_enable = "ena0";
defparam ram_block1a56.clk0_input_clock_enable = "ena0";
defparam ram_block1a56.clk1_core_clock_enable = "ena1";
defparam ram_block1a56.clk1_input_clock_enable = "ena1";
defparam ram_block1a56.data_interleave_offset_in_bits = 1;
defparam ram_block1a56.data_interleave_width_in_bits = 1;
defparam ram_block1a56.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a56.init_file_layout = "port_a";
defparam ram_block1a56.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a56.operation_mode = "bidir_dual_port";
defparam ram_block1a56.port_a_address_clear = "none";
defparam ram_block1a56.port_a_address_width = 13;
defparam ram_block1a56.port_a_byte_enable_mask_width = 1;
defparam ram_block1a56.port_a_byte_size = 1;
defparam ram_block1a56.port_a_data_out_clear = "none";
defparam ram_block1a56.port_a_data_out_clock = "none";
defparam ram_block1a56.port_a_data_width = 1;
defparam ram_block1a56.port_a_first_address = 0;
defparam ram_block1a56.port_a_first_bit_number = 56;
defparam ram_block1a56.port_a_last_address = 8191;
defparam ram_block1a56.port_a_logical_ram_depth = 16384;
defparam ram_block1a56.port_a_logical_ram_width = 64;
defparam ram_block1a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a56.port_b_address_clear = "none";
defparam ram_block1a56.port_b_address_clock = "clock1";
defparam ram_block1a56.port_b_address_width = 13;
defparam ram_block1a56.port_b_byte_enable_clock = "clock1";
defparam ram_block1a56.port_b_byte_enable_mask_width = 1;
defparam ram_block1a56.port_b_byte_size = 1;
defparam ram_block1a56.port_b_data_in_clock = "clock1";
defparam ram_block1a56.port_b_data_out_clear = "none";
defparam ram_block1a56.port_b_data_out_clock = "none";
defparam ram_block1a56.port_b_data_width = 1;
defparam ram_block1a56.port_b_first_address = 0;
defparam ram_block1a56.port_b_first_bit_number = 56;
defparam ram_block1a56.port_b_last_address = 8191;
defparam ram_block1a56.port_b_logical_ram_depth = 16384;
defparam ram_block1a56.port_b_logical_ram_width = 64;
defparam ram_block1a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a56.port_b_read_enable_clock = "clock1";
defparam ram_block1a56.port_b_write_enable_clock = "clock1";
defparam ram_block1a56.ram_block_type = "auto";
defparam ram_block1a56.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a56.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a56.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a56.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a121(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[57]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[57]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a121_PORTADATAOUT_bus),
	.portbdataout(ram_block1a121_PORTBDATAOUT_bus));
defparam ram_block1a121.clk0_core_clock_enable = "ena0";
defparam ram_block1a121.clk0_input_clock_enable = "ena0";
defparam ram_block1a121.clk1_core_clock_enable = "ena1";
defparam ram_block1a121.clk1_input_clock_enable = "ena1";
defparam ram_block1a121.data_interleave_offset_in_bits = 1;
defparam ram_block1a121.data_interleave_width_in_bits = 1;
defparam ram_block1a121.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a121.init_file_layout = "port_a";
defparam ram_block1a121.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a121.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a121.operation_mode = "bidir_dual_port";
defparam ram_block1a121.port_a_address_clear = "none";
defparam ram_block1a121.port_a_address_width = 13;
defparam ram_block1a121.port_a_byte_enable_mask_width = 1;
defparam ram_block1a121.port_a_byte_size = 1;
defparam ram_block1a121.port_a_data_out_clear = "none";
defparam ram_block1a121.port_a_data_out_clock = "none";
defparam ram_block1a121.port_a_data_width = 1;
defparam ram_block1a121.port_a_first_address = 8192;
defparam ram_block1a121.port_a_first_bit_number = 57;
defparam ram_block1a121.port_a_last_address = 16383;
defparam ram_block1a121.port_a_logical_ram_depth = 16384;
defparam ram_block1a121.port_a_logical_ram_width = 64;
defparam ram_block1a121.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a121.port_b_address_clear = "none";
defparam ram_block1a121.port_b_address_clock = "clock1";
defparam ram_block1a121.port_b_address_width = 13;
defparam ram_block1a121.port_b_byte_enable_clock = "clock1";
defparam ram_block1a121.port_b_byte_enable_mask_width = 1;
defparam ram_block1a121.port_b_byte_size = 1;
defparam ram_block1a121.port_b_data_in_clock = "clock1";
defparam ram_block1a121.port_b_data_out_clear = "none";
defparam ram_block1a121.port_b_data_out_clock = "none";
defparam ram_block1a121.port_b_data_width = 1;
defparam ram_block1a121.port_b_first_address = 8192;
defparam ram_block1a121.port_b_first_bit_number = 57;
defparam ram_block1a121.port_b_last_address = 16383;
defparam ram_block1a121.port_b_logical_ram_depth = 16384;
defparam ram_block1a121.port_b_logical_ram_width = 64;
defparam ram_block1a121.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a121.port_b_read_enable_clock = "clock1";
defparam ram_block1a121.port_b_write_enable_clock = "clock1";
defparam ram_block1a121.ram_block_type = "auto";
defparam ram_block1a121.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a121.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a121.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a121.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a57(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[57]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[57]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a57_PORTADATAOUT_bus),
	.portbdataout(ram_block1a57_PORTBDATAOUT_bus));
defparam ram_block1a57.clk0_core_clock_enable = "ena0";
defparam ram_block1a57.clk0_input_clock_enable = "ena0";
defparam ram_block1a57.clk1_core_clock_enable = "ena1";
defparam ram_block1a57.clk1_input_clock_enable = "ena1";
defparam ram_block1a57.data_interleave_offset_in_bits = 1;
defparam ram_block1a57.data_interleave_width_in_bits = 1;
defparam ram_block1a57.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a57.init_file_layout = "port_a";
defparam ram_block1a57.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a57.operation_mode = "bidir_dual_port";
defparam ram_block1a57.port_a_address_clear = "none";
defparam ram_block1a57.port_a_address_width = 13;
defparam ram_block1a57.port_a_byte_enable_mask_width = 1;
defparam ram_block1a57.port_a_byte_size = 1;
defparam ram_block1a57.port_a_data_out_clear = "none";
defparam ram_block1a57.port_a_data_out_clock = "none";
defparam ram_block1a57.port_a_data_width = 1;
defparam ram_block1a57.port_a_first_address = 0;
defparam ram_block1a57.port_a_first_bit_number = 57;
defparam ram_block1a57.port_a_last_address = 8191;
defparam ram_block1a57.port_a_logical_ram_depth = 16384;
defparam ram_block1a57.port_a_logical_ram_width = 64;
defparam ram_block1a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a57.port_b_address_clear = "none";
defparam ram_block1a57.port_b_address_clock = "clock1";
defparam ram_block1a57.port_b_address_width = 13;
defparam ram_block1a57.port_b_byte_enable_clock = "clock1";
defparam ram_block1a57.port_b_byte_enable_mask_width = 1;
defparam ram_block1a57.port_b_byte_size = 1;
defparam ram_block1a57.port_b_data_in_clock = "clock1";
defparam ram_block1a57.port_b_data_out_clear = "none";
defparam ram_block1a57.port_b_data_out_clock = "none";
defparam ram_block1a57.port_b_data_width = 1;
defparam ram_block1a57.port_b_first_address = 0;
defparam ram_block1a57.port_b_first_bit_number = 57;
defparam ram_block1a57.port_b_last_address = 8191;
defparam ram_block1a57.port_b_logical_ram_depth = 16384;
defparam ram_block1a57.port_b_logical_ram_width = 64;
defparam ram_block1a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a57.port_b_read_enable_clock = "clock1";
defparam ram_block1a57.port_b_write_enable_clock = "clock1";
defparam ram_block1a57.ram_block_type = "auto";
defparam ram_block1a57.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a57.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a57.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a57.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a122(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[58]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[58]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a122_PORTADATAOUT_bus),
	.portbdataout(ram_block1a122_PORTBDATAOUT_bus));
defparam ram_block1a122.clk0_core_clock_enable = "ena0";
defparam ram_block1a122.clk0_input_clock_enable = "ena0";
defparam ram_block1a122.clk1_core_clock_enable = "ena1";
defparam ram_block1a122.clk1_input_clock_enable = "ena1";
defparam ram_block1a122.data_interleave_offset_in_bits = 1;
defparam ram_block1a122.data_interleave_width_in_bits = 1;
defparam ram_block1a122.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a122.init_file_layout = "port_a";
defparam ram_block1a122.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a122.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a122.operation_mode = "bidir_dual_port";
defparam ram_block1a122.port_a_address_clear = "none";
defparam ram_block1a122.port_a_address_width = 13;
defparam ram_block1a122.port_a_byte_enable_mask_width = 1;
defparam ram_block1a122.port_a_byte_size = 1;
defparam ram_block1a122.port_a_data_out_clear = "none";
defparam ram_block1a122.port_a_data_out_clock = "none";
defparam ram_block1a122.port_a_data_width = 1;
defparam ram_block1a122.port_a_first_address = 8192;
defparam ram_block1a122.port_a_first_bit_number = 58;
defparam ram_block1a122.port_a_last_address = 16383;
defparam ram_block1a122.port_a_logical_ram_depth = 16384;
defparam ram_block1a122.port_a_logical_ram_width = 64;
defparam ram_block1a122.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a122.port_b_address_clear = "none";
defparam ram_block1a122.port_b_address_clock = "clock1";
defparam ram_block1a122.port_b_address_width = 13;
defparam ram_block1a122.port_b_byte_enable_clock = "clock1";
defparam ram_block1a122.port_b_byte_enable_mask_width = 1;
defparam ram_block1a122.port_b_byte_size = 1;
defparam ram_block1a122.port_b_data_in_clock = "clock1";
defparam ram_block1a122.port_b_data_out_clear = "none";
defparam ram_block1a122.port_b_data_out_clock = "none";
defparam ram_block1a122.port_b_data_width = 1;
defparam ram_block1a122.port_b_first_address = 8192;
defparam ram_block1a122.port_b_first_bit_number = 58;
defparam ram_block1a122.port_b_last_address = 16383;
defparam ram_block1a122.port_b_logical_ram_depth = 16384;
defparam ram_block1a122.port_b_logical_ram_width = 64;
defparam ram_block1a122.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a122.port_b_read_enable_clock = "clock1";
defparam ram_block1a122.port_b_write_enable_clock = "clock1";
defparam ram_block1a122.ram_block_type = "auto";
defparam ram_block1a122.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a122.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a122.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a122.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a58(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[58]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[58]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a58_PORTADATAOUT_bus),
	.portbdataout(ram_block1a58_PORTBDATAOUT_bus));
defparam ram_block1a58.clk0_core_clock_enable = "ena0";
defparam ram_block1a58.clk0_input_clock_enable = "ena0";
defparam ram_block1a58.clk1_core_clock_enable = "ena1";
defparam ram_block1a58.clk1_input_clock_enable = "ena1";
defparam ram_block1a58.data_interleave_offset_in_bits = 1;
defparam ram_block1a58.data_interleave_width_in_bits = 1;
defparam ram_block1a58.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a58.init_file_layout = "port_a";
defparam ram_block1a58.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a58.operation_mode = "bidir_dual_port";
defparam ram_block1a58.port_a_address_clear = "none";
defparam ram_block1a58.port_a_address_width = 13;
defparam ram_block1a58.port_a_byte_enable_mask_width = 1;
defparam ram_block1a58.port_a_byte_size = 1;
defparam ram_block1a58.port_a_data_out_clear = "none";
defparam ram_block1a58.port_a_data_out_clock = "none";
defparam ram_block1a58.port_a_data_width = 1;
defparam ram_block1a58.port_a_first_address = 0;
defparam ram_block1a58.port_a_first_bit_number = 58;
defparam ram_block1a58.port_a_last_address = 8191;
defparam ram_block1a58.port_a_logical_ram_depth = 16384;
defparam ram_block1a58.port_a_logical_ram_width = 64;
defparam ram_block1a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a58.port_b_address_clear = "none";
defparam ram_block1a58.port_b_address_clock = "clock1";
defparam ram_block1a58.port_b_address_width = 13;
defparam ram_block1a58.port_b_byte_enable_clock = "clock1";
defparam ram_block1a58.port_b_byte_enable_mask_width = 1;
defparam ram_block1a58.port_b_byte_size = 1;
defparam ram_block1a58.port_b_data_in_clock = "clock1";
defparam ram_block1a58.port_b_data_out_clear = "none";
defparam ram_block1a58.port_b_data_out_clock = "none";
defparam ram_block1a58.port_b_data_width = 1;
defparam ram_block1a58.port_b_first_address = 0;
defparam ram_block1a58.port_b_first_bit_number = 58;
defparam ram_block1a58.port_b_last_address = 8191;
defparam ram_block1a58.port_b_logical_ram_depth = 16384;
defparam ram_block1a58.port_b_logical_ram_width = 64;
defparam ram_block1a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a58.port_b_read_enable_clock = "clock1";
defparam ram_block1a58.port_b_write_enable_clock = "clock1";
defparam ram_block1a58.ram_block_type = "auto";
defparam ram_block1a58.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a58.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a58.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a58.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a123(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[59]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[59]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a123_PORTADATAOUT_bus),
	.portbdataout(ram_block1a123_PORTBDATAOUT_bus));
defparam ram_block1a123.clk0_core_clock_enable = "ena0";
defparam ram_block1a123.clk0_input_clock_enable = "ena0";
defparam ram_block1a123.clk1_core_clock_enable = "ena1";
defparam ram_block1a123.clk1_input_clock_enable = "ena1";
defparam ram_block1a123.data_interleave_offset_in_bits = 1;
defparam ram_block1a123.data_interleave_width_in_bits = 1;
defparam ram_block1a123.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a123.init_file_layout = "port_a";
defparam ram_block1a123.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a123.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a123.operation_mode = "bidir_dual_port";
defparam ram_block1a123.port_a_address_clear = "none";
defparam ram_block1a123.port_a_address_width = 13;
defparam ram_block1a123.port_a_byte_enable_mask_width = 1;
defparam ram_block1a123.port_a_byte_size = 1;
defparam ram_block1a123.port_a_data_out_clear = "none";
defparam ram_block1a123.port_a_data_out_clock = "none";
defparam ram_block1a123.port_a_data_width = 1;
defparam ram_block1a123.port_a_first_address = 8192;
defparam ram_block1a123.port_a_first_bit_number = 59;
defparam ram_block1a123.port_a_last_address = 16383;
defparam ram_block1a123.port_a_logical_ram_depth = 16384;
defparam ram_block1a123.port_a_logical_ram_width = 64;
defparam ram_block1a123.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a123.port_b_address_clear = "none";
defparam ram_block1a123.port_b_address_clock = "clock1";
defparam ram_block1a123.port_b_address_width = 13;
defparam ram_block1a123.port_b_byte_enable_clock = "clock1";
defparam ram_block1a123.port_b_byte_enable_mask_width = 1;
defparam ram_block1a123.port_b_byte_size = 1;
defparam ram_block1a123.port_b_data_in_clock = "clock1";
defparam ram_block1a123.port_b_data_out_clear = "none";
defparam ram_block1a123.port_b_data_out_clock = "none";
defparam ram_block1a123.port_b_data_width = 1;
defparam ram_block1a123.port_b_first_address = 8192;
defparam ram_block1a123.port_b_first_bit_number = 59;
defparam ram_block1a123.port_b_last_address = 16383;
defparam ram_block1a123.port_b_logical_ram_depth = 16384;
defparam ram_block1a123.port_b_logical_ram_width = 64;
defparam ram_block1a123.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a123.port_b_read_enable_clock = "clock1";
defparam ram_block1a123.port_b_write_enable_clock = "clock1";
defparam ram_block1a123.ram_block_type = "auto";
defparam ram_block1a123.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a123.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a123.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a123.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a59(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[59]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[59]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a59_PORTADATAOUT_bus),
	.portbdataout(ram_block1a59_PORTBDATAOUT_bus));
defparam ram_block1a59.clk0_core_clock_enable = "ena0";
defparam ram_block1a59.clk0_input_clock_enable = "ena0";
defparam ram_block1a59.clk1_core_clock_enable = "ena1";
defparam ram_block1a59.clk1_input_clock_enable = "ena1";
defparam ram_block1a59.data_interleave_offset_in_bits = 1;
defparam ram_block1a59.data_interleave_width_in_bits = 1;
defparam ram_block1a59.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a59.init_file_layout = "port_a";
defparam ram_block1a59.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a59.operation_mode = "bidir_dual_port";
defparam ram_block1a59.port_a_address_clear = "none";
defparam ram_block1a59.port_a_address_width = 13;
defparam ram_block1a59.port_a_byte_enable_mask_width = 1;
defparam ram_block1a59.port_a_byte_size = 1;
defparam ram_block1a59.port_a_data_out_clear = "none";
defparam ram_block1a59.port_a_data_out_clock = "none";
defparam ram_block1a59.port_a_data_width = 1;
defparam ram_block1a59.port_a_first_address = 0;
defparam ram_block1a59.port_a_first_bit_number = 59;
defparam ram_block1a59.port_a_last_address = 8191;
defparam ram_block1a59.port_a_logical_ram_depth = 16384;
defparam ram_block1a59.port_a_logical_ram_width = 64;
defparam ram_block1a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a59.port_b_address_clear = "none";
defparam ram_block1a59.port_b_address_clock = "clock1";
defparam ram_block1a59.port_b_address_width = 13;
defparam ram_block1a59.port_b_byte_enable_clock = "clock1";
defparam ram_block1a59.port_b_byte_enable_mask_width = 1;
defparam ram_block1a59.port_b_byte_size = 1;
defparam ram_block1a59.port_b_data_in_clock = "clock1";
defparam ram_block1a59.port_b_data_out_clear = "none";
defparam ram_block1a59.port_b_data_out_clock = "none";
defparam ram_block1a59.port_b_data_width = 1;
defparam ram_block1a59.port_b_first_address = 0;
defparam ram_block1a59.port_b_first_bit_number = 59;
defparam ram_block1a59.port_b_last_address = 8191;
defparam ram_block1a59.port_b_logical_ram_depth = 16384;
defparam ram_block1a59.port_b_logical_ram_width = 64;
defparam ram_block1a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a59.port_b_read_enable_clock = "clock1";
defparam ram_block1a59.port_b_write_enable_clock = "clock1";
defparam ram_block1a59.ram_block_type = "auto";
defparam ram_block1a59.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a59.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a59.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a59.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a124(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[60]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[60]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a124_PORTADATAOUT_bus),
	.portbdataout(ram_block1a124_PORTBDATAOUT_bus));
defparam ram_block1a124.clk0_core_clock_enable = "ena0";
defparam ram_block1a124.clk0_input_clock_enable = "ena0";
defparam ram_block1a124.clk1_core_clock_enable = "ena1";
defparam ram_block1a124.clk1_input_clock_enable = "ena1";
defparam ram_block1a124.data_interleave_offset_in_bits = 1;
defparam ram_block1a124.data_interleave_width_in_bits = 1;
defparam ram_block1a124.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a124.init_file_layout = "port_a";
defparam ram_block1a124.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a124.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a124.operation_mode = "bidir_dual_port";
defparam ram_block1a124.port_a_address_clear = "none";
defparam ram_block1a124.port_a_address_width = 13;
defparam ram_block1a124.port_a_byte_enable_mask_width = 1;
defparam ram_block1a124.port_a_byte_size = 1;
defparam ram_block1a124.port_a_data_out_clear = "none";
defparam ram_block1a124.port_a_data_out_clock = "none";
defparam ram_block1a124.port_a_data_width = 1;
defparam ram_block1a124.port_a_first_address = 8192;
defparam ram_block1a124.port_a_first_bit_number = 60;
defparam ram_block1a124.port_a_last_address = 16383;
defparam ram_block1a124.port_a_logical_ram_depth = 16384;
defparam ram_block1a124.port_a_logical_ram_width = 64;
defparam ram_block1a124.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a124.port_b_address_clear = "none";
defparam ram_block1a124.port_b_address_clock = "clock1";
defparam ram_block1a124.port_b_address_width = 13;
defparam ram_block1a124.port_b_byte_enable_clock = "clock1";
defparam ram_block1a124.port_b_byte_enable_mask_width = 1;
defparam ram_block1a124.port_b_byte_size = 1;
defparam ram_block1a124.port_b_data_in_clock = "clock1";
defparam ram_block1a124.port_b_data_out_clear = "none";
defparam ram_block1a124.port_b_data_out_clock = "none";
defparam ram_block1a124.port_b_data_width = 1;
defparam ram_block1a124.port_b_first_address = 8192;
defparam ram_block1a124.port_b_first_bit_number = 60;
defparam ram_block1a124.port_b_last_address = 16383;
defparam ram_block1a124.port_b_logical_ram_depth = 16384;
defparam ram_block1a124.port_b_logical_ram_width = 64;
defparam ram_block1a124.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a124.port_b_read_enable_clock = "clock1";
defparam ram_block1a124.port_b_write_enable_clock = "clock1";
defparam ram_block1a124.ram_block_type = "auto";
defparam ram_block1a124.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a124.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a124.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a124.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a60(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[60]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[60]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a60_PORTADATAOUT_bus),
	.portbdataout(ram_block1a60_PORTBDATAOUT_bus));
defparam ram_block1a60.clk0_core_clock_enable = "ena0";
defparam ram_block1a60.clk0_input_clock_enable = "ena0";
defparam ram_block1a60.clk1_core_clock_enable = "ena1";
defparam ram_block1a60.clk1_input_clock_enable = "ena1";
defparam ram_block1a60.data_interleave_offset_in_bits = 1;
defparam ram_block1a60.data_interleave_width_in_bits = 1;
defparam ram_block1a60.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a60.init_file_layout = "port_a";
defparam ram_block1a60.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a60.operation_mode = "bidir_dual_port";
defparam ram_block1a60.port_a_address_clear = "none";
defparam ram_block1a60.port_a_address_width = 13;
defparam ram_block1a60.port_a_byte_enable_mask_width = 1;
defparam ram_block1a60.port_a_byte_size = 1;
defparam ram_block1a60.port_a_data_out_clear = "none";
defparam ram_block1a60.port_a_data_out_clock = "none";
defparam ram_block1a60.port_a_data_width = 1;
defparam ram_block1a60.port_a_first_address = 0;
defparam ram_block1a60.port_a_first_bit_number = 60;
defparam ram_block1a60.port_a_last_address = 8191;
defparam ram_block1a60.port_a_logical_ram_depth = 16384;
defparam ram_block1a60.port_a_logical_ram_width = 64;
defparam ram_block1a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a60.port_b_address_clear = "none";
defparam ram_block1a60.port_b_address_clock = "clock1";
defparam ram_block1a60.port_b_address_width = 13;
defparam ram_block1a60.port_b_byte_enable_clock = "clock1";
defparam ram_block1a60.port_b_byte_enable_mask_width = 1;
defparam ram_block1a60.port_b_byte_size = 1;
defparam ram_block1a60.port_b_data_in_clock = "clock1";
defparam ram_block1a60.port_b_data_out_clear = "none";
defparam ram_block1a60.port_b_data_out_clock = "none";
defparam ram_block1a60.port_b_data_width = 1;
defparam ram_block1a60.port_b_first_address = 0;
defparam ram_block1a60.port_b_first_bit_number = 60;
defparam ram_block1a60.port_b_last_address = 8191;
defparam ram_block1a60.port_b_logical_ram_depth = 16384;
defparam ram_block1a60.port_b_logical_ram_width = 64;
defparam ram_block1a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a60.port_b_read_enable_clock = "clock1";
defparam ram_block1a60.port_b_write_enable_clock = "clock1";
defparam ram_block1a60.ram_block_type = "auto";
defparam ram_block1a60.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a60.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a60.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a60.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a125(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[61]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[61]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a125_PORTADATAOUT_bus),
	.portbdataout(ram_block1a125_PORTBDATAOUT_bus));
defparam ram_block1a125.clk0_core_clock_enable = "ena0";
defparam ram_block1a125.clk0_input_clock_enable = "ena0";
defparam ram_block1a125.clk1_core_clock_enable = "ena1";
defparam ram_block1a125.clk1_input_clock_enable = "ena1";
defparam ram_block1a125.data_interleave_offset_in_bits = 1;
defparam ram_block1a125.data_interleave_width_in_bits = 1;
defparam ram_block1a125.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a125.init_file_layout = "port_a";
defparam ram_block1a125.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a125.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a125.operation_mode = "bidir_dual_port";
defparam ram_block1a125.port_a_address_clear = "none";
defparam ram_block1a125.port_a_address_width = 13;
defparam ram_block1a125.port_a_byte_enable_mask_width = 1;
defparam ram_block1a125.port_a_byte_size = 1;
defparam ram_block1a125.port_a_data_out_clear = "none";
defparam ram_block1a125.port_a_data_out_clock = "none";
defparam ram_block1a125.port_a_data_width = 1;
defparam ram_block1a125.port_a_first_address = 8192;
defparam ram_block1a125.port_a_first_bit_number = 61;
defparam ram_block1a125.port_a_last_address = 16383;
defparam ram_block1a125.port_a_logical_ram_depth = 16384;
defparam ram_block1a125.port_a_logical_ram_width = 64;
defparam ram_block1a125.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a125.port_b_address_clear = "none";
defparam ram_block1a125.port_b_address_clock = "clock1";
defparam ram_block1a125.port_b_address_width = 13;
defparam ram_block1a125.port_b_byte_enable_clock = "clock1";
defparam ram_block1a125.port_b_byte_enable_mask_width = 1;
defparam ram_block1a125.port_b_byte_size = 1;
defparam ram_block1a125.port_b_data_in_clock = "clock1";
defparam ram_block1a125.port_b_data_out_clear = "none";
defparam ram_block1a125.port_b_data_out_clock = "none";
defparam ram_block1a125.port_b_data_width = 1;
defparam ram_block1a125.port_b_first_address = 8192;
defparam ram_block1a125.port_b_first_bit_number = 61;
defparam ram_block1a125.port_b_last_address = 16383;
defparam ram_block1a125.port_b_logical_ram_depth = 16384;
defparam ram_block1a125.port_b_logical_ram_width = 64;
defparam ram_block1a125.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a125.port_b_read_enable_clock = "clock1";
defparam ram_block1a125.port_b_write_enable_clock = "clock1";
defparam ram_block1a125.ram_block_type = "auto";
defparam ram_block1a125.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a125.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a125.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a125.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a61(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[61]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[61]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a61_PORTADATAOUT_bus),
	.portbdataout(ram_block1a61_PORTBDATAOUT_bus));
defparam ram_block1a61.clk0_core_clock_enable = "ena0";
defparam ram_block1a61.clk0_input_clock_enable = "ena0";
defparam ram_block1a61.clk1_core_clock_enable = "ena1";
defparam ram_block1a61.clk1_input_clock_enable = "ena1";
defparam ram_block1a61.data_interleave_offset_in_bits = 1;
defparam ram_block1a61.data_interleave_width_in_bits = 1;
defparam ram_block1a61.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a61.init_file_layout = "port_a";
defparam ram_block1a61.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a61.operation_mode = "bidir_dual_port";
defparam ram_block1a61.port_a_address_clear = "none";
defparam ram_block1a61.port_a_address_width = 13;
defparam ram_block1a61.port_a_byte_enable_mask_width = 1;
defparam ram_block1a61.port_a_byte_size = 1;
defparam ram_block1a61.port_a_data_out_clear = "none";
defparam ram_block1a61.port_a_data_out_clock = "none";
defparam ram_block1a61.port_a_data_width = 1;
defparam ram_block1a61.port_a_first_address = 0;
defparam ram_block1a61.port_a_first_bit_number = 61;
defparam ram_block1a61.port_a_last_address = 8191;
defparam ram_block1a61.port_a_logical_ram_depth = 16384;
defparam ram_block1a61.port_a_logical_ram_width = 64;
defparam ram_block1a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a61.port_b_address_clear = "none";
defparam ram_block1a61.port_b_address_clock = "clock1";
defparam ram_block1a61.port_b_address_width = 13;
defparam ram_block1a61.port_b_byte_enable_clock = "clock1";
defparam ram_block1a61.port_b_byte_enable_mask_width = 1;
defparam ram_block1a61.port_b_byte_size = 1;
defparam ram_block1a61.port_b_data_in_clock = "clock1";
defparam ram_block1a61.port_b_data_out_clear = "none";
defparam ram_block1a61.port_b_data_out_clock = "none";
defparam ram_block1a61.port_b_data_width = 1;
defparam ram_block1a61.port_b_first_address = 0;
defparam ram_block1a61.port_b_first_bit_number = 61;
defparam ram_block1a61.port_b_last_address = 8191;
defparam ram_block1a61.port_b_logical_ram_depth = 16384;
defparam ram_block1a61.port_b_logical_ram_width = 64;
defparam ram_block1a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a61.port_b_read_enable_clock = "clock1";
defparam ram_block1a61.port_b_write_enable_clock = "clock1";
defparam ram_block1a61.ram_block_type = "auto";
defparam ram_block1a61.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a61.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a61.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a61.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a126(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[62]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[62]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a126_PORTADATAOUT_bus),
	.portbdataout(ram_block1a126_PORTBDATAOUT_bus));
defparam ram_block1a126.clk0_core_clock_enable = "ena0";
defparam ram_block1a126.clk0_input_clock_enable = "ena0";
defparam ram_block1a126.clk1_core_clock_enable = "ena1";
defparam ram_block1a126.clk1_input_clock_enable = "ena1";
defparam ram_block1a126.data_interleave_offset_in_bits = 1;
defparam ram_block1a126.data_interleave_width_in_bits = 1;
defparam ram_block1a126.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a126.init_file_layout = "port_a";
defparam ram_block1a126.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a126.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a126.operation_mode = "bidir_dual_port";
defparam ram_block1a126.port_a_address_clear = "none";
defparam ram_block1a126.port_a_address_width = 13;
defparam ram_block1a126.port_a_byte_enable_mask_width = 1;
defparam ram_block1a126.port_a_byte_size = 1;
defparam ram_block1a126.port_a_data_out_clear = "none";
defparam ram_block1a126.port_a_data_out_clock = "none";
defparam ram_block1a126.port_a_data_width = 1;
defparam ram_block1a126.port_a_first_address = 8192;
defparam ram_block1a126.port_a_first_bit_number = 62;
defparam ram_block1a126.port_a_last_address = 16383;
defparam ram_block1a126.port_a_logical_ram_depth = 16384;
defparam ram_block1a126.port_a_logical_ram_width = 64;
defparam ram_block1a126.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a126.port_b_address_clear = "none";
defparam ram_block1a126.port_b_address_clock = "clock1";
defparam ram_block1a126.port_b_address_width = 13;
defparam ram_block1a126.port_b_byte_enable_clock = "clock1";
defparam ram_block1a126.port_b_byte_enable_mask_width = 1;
defparam ram_block1a126.port_b_byte_size = 1;
defparam ram_block1a126.port_b_data_in_clock = "clock1";
defparam ram_block1a126.port_b_data_out_clear = "none";
defparam ram_block1a126.port_b_data_out_clock = "none";
defparam ram_block1a126.port_b_data_width = 1;
defparam ram_block1a126.port_b_first_address = 8192;
defparam ram_block1a126.port_b_first_bit_number = 62;
defparam ram_block1a126.port_b_last_address = 16383;
defparam ram_block1a126.port_b_logical_ram_depth = 16384;
defparam ram_block1a126.port_b_logical_ram_width = 64;
defparam ram_block1a126.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a126.port_b_read_enable_clock = "clock1";
defparam ram_block1a126.port_b_write_enable_clock = "clock1";
defparam ram_block1a126.ram_block_type = "auto";
defparam ram_block1a126.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a126.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a126.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a126.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a62(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[62]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[62]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a62_PORTADATAOUT_bus),
	.portbdataout(ram_block1a62_PORTBDATAOUT_bus));
defparam ram_block1a62.clk0_core_clock_enable = "ena0";
defparam ram_block1a62.clk0_input_clock_enable = "ena0";
defparam ram_block1a62.clk1_core_clock_enable = "ena1";
defparam ram_block1a62.clk1_input_clock_enable = "ena1";
defparam ram_block1a62.data_interleave_offset_in_bits = 1;
defparam ram_block1a62.data_interleave_width_in_bits = 1;
defparam ram_block1a62.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a62.init_file_layout = "port_a";
defparam ram_block1a62.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a62.operation_mode = "bidir_dual_port";
defparam ram_block1a62.port_a_address_clear = "none";
defparam ram_block1a62.port_a_address_width = 13;
defparam ram_block1a62.port_a_byte_enable_mask_width = 1;
defparam ram_block1a62.port_a_byte_size = 1;
defparam ram_block1a62.port_a_data_out_clear = "none";
defparam ram_block1a62.port_a_data_out_clock = "none";
defparam ram_block1a62.port_a_data_width = 1;
defparam ram_block1a62.port_a_first_address = 0;
defparam ram_block1a62.port_a_first_bit_number = 62;
defparam ram_block1a62.port_a_last_address = 8191;
defparam ram_block1a62.port_a_logical_ram_depth = 16384;
defparam ram_block1a62.port_a_logical_ram_width = 64;
defparam ram_block1a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a62.port_b_address_clear = "none";
defparam ram_block1a62.port_b_address_clock = "clock1";
defparam ram_block1a62.port_b_address_width = 13;
defparam ram_block1a62.port_b_byte_enable_clock = "clock1";
defparam ram_block1a62.port_b_byte_enable_mask_width = 1;
defparam ram_block1a62.port_b_byte_size = 1;
defparam ram_block1a62.port_b_data_in_clock = "clock1";
defparam ram_block1a62.port_b_data_out_clear = "none";
defparam ram_block1a62.port_b_data_out_clock = "none";
defparam ram_block1a62.port_b_data_width = 1;
defparam ram_block1a62.port_b_first_address = 0;
defparam ram_block1a62.port_b_first_bit_number = 62;
defparam ram_block1a62.port_b_last_address = 8191;
defparam ram_block1a62.port_b_logical_ram_depth = 16384;
defparam ram_block1a62.port_b_logical_ram_width = 64;
defparam ram_block1a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a62.port_b_read_enable_clock = "clock1";
defparam ram_block1a62.port_b_write_enable_clock = "clock1";
defparam ram_block1a62.ram_block_type = "auto";
defparam ram_block1a62.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a62.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a62.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a62.mem_init0 = 2048'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

cycloneiv_ram_block ram_block1a127(
	.portawe(\decode2|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[63]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[63]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a127_PORTADATAOUT_bus),
	.portbdataout(ram_block1a127_PORTBDATAOUT_bus));
defparam ram_block1a127.clk0_core_clock_enable = "ena0";
defparam ram_block1a127.clk0_input_clock_enable = "ena0";
defparam ram_block1a127.clk1_core_clock_enable = "ena1";
defparam ram_block1a127.clk1_input_clock_enable = "ena1";
defparam ram_block1a127.data_interleave_offset_in_bits = 1;
defparam ram_block1a127.data_interleave_width_in_bits = 1;
defparam ram_block1a127.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a127.init_file_layout = "port_a";
defparam ram_block1a127.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a127.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a127.operation_mode = "bidir_dual_port";
defparam ram_block1a127.port_a_address_clear = "none";
defparam ram_block1a127.port_a_address_width = 13;
defparam ram_block1a127.port_a_byte_enable_mask_width = 1;
defparam ram_block1a127.port_a_byte_size = 1;
defparam ram_block1a127.port_a_data_out_clear = "none";
defparam ram_block1a127.port_a_data_out_clock = "none";
defparam ram_block1a127.port_a_data_width = 1;
defparam ram_block1a127.port_a_first_address = 8192;
defparam ram_block1a127.port_a_first_bit_number = 63;
defparam ram_block1a127.port_a_last_address = 16383;
defparam ram_block1a127.port_a_logical_ram_depth = 16384;
defparam ram_block1a127.port_a_logical_ram_width = 64;
defparam ram_block1a127.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a127.port_b_address_clear = "none";
defparam ram_block1a127.port_b_address_clock = "clock1";
defparam ram_block1a127.port_b_address_width = 13;
defparam ram_block1a127.port_b_byte_enable_clock = "clock1";
defparam ram_block1a127.port_b_byte_enable_mask_width = 1;
defparam ram_block1a127.port_b_byte_size = 1;
defparam ram_block1a127.port_b_data_in_clock = "clock1";
defparam ram_block1a127.port_b_data_out_clear = "none";
defparam ram_block1a127.port_b_data_out_clock = "none";
defparam ram_block1a127.port_b_data_width = 1;
defparam ram_block1a127.port_b_first_address = 8192;
defparam ram_block1a127.port_b_first_bit_number = 63;
defparam ram_block1a127.port_b_last_address = 16383;
defparam ram_block1a127.port_b_logical_ram_depth = 16384;
defparam ram_block1a127.port_b_logical_ram_width = 64;
defparam ram_block1a127.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a127.port_b_read_enable_clock = "clock1";
defparam ram_block1a127.port_b_write_enable_clock = "clock1";
defparam ram_block1a127.ram_block_type = "auto";
defparam ram_block1a127.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a127.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a127.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a127.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

cycloneiv_ram_block ram_block1a63(
	.portawe(\decode2|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode3|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock1),
	.clk1(clock1),
	.ena0(clocken0),
	.ena1(clocken1),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[63]}),
	.portaaddr({gnd,gnd,gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[7]}),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_b[63]}),
	.portbaddr({gnd,gnd,gnd,address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_b[7]}),
	.portadataout(ram_block1a63_PORTADATAOUT_bus),
	.portbdataout(ram_block1a63_PORTBDATAOUT_bus));
defparam ram_block1a63.clk0_core_clock_enable = "ena0";
defparam ram_block1a63.clk0_input_clock_enable = "ena0";
defparam ram_block1a63.clk1_core_clock_enable = "ena1";
defparam ram_block1a63.clk1_input_clock_enable = "ena1";
defparam ram_block1a63.data_interleave_offset_in_bits = 1;
defparam ram_block1a63.data_interleave_width_in_bits = 1;
defparam ram_block1a63.init_file = "D:/Cinna-BoN-FPGA/qtest/qtest.hex";
defparam ram_block1a63.init_file_layout = "port_a";
defparam ram_block1a63.logical_ram_name = "qtestpd_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_6342:auto_generated|ALTSYNCRAM";
defparam ram_block1a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a63.operation_mode = "bidir_dual_port";
defparam ram_block1a63.port_a_address_clear = "none";
defparam ram_block1a63.port_a_address_width = 13;
defparam ram_block1a63.port_a_byte_enable_mask_width = 1;
defparam ram_block1a63.port_a_byte_size = 1;
defparam ram_block1a63.port_a_data_out_clear = "none";
defparam ram_block1a63.port_a_data_out_clock = "none";
defparam ram_block1a63.port_a_data_width = 1;
defparam ram_block1a63.port_a_first_address = 0;
defparam ram_block1a63.port_a_first_bit_number = 63;
defparam ram_block1a63.port_a_last_address = 8191;
defparam ram_block1a63.port_a_logical_ram_depth = 16384;
defparam ram_block1a63.port_a_logical_ram_width = 64;
defparam ram_block1a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a63.port_b_address_clear = "none";
defparam ram_block1a63.port_b_address_clock = "clock1";
defparam ram_block1a63.port_b_address_width = 13;
defparam ram_block1a63.port_b_byte_enable_clock = "clock1";
defparam ram_block1a63.port_b_byte_enable_mask_width = 1;
defparam ram_block1a63.port_b_byte_size = 1;
defparam ram_block1a63.port_b_data_in_clock = "clock1";
defparam ram_block1a63.port_b_data_out_clear = "none";
defparam ram_block1a63.port_b_data_out_clock = "none";
defparam ram_block1a63.port_b_data_width = 1;
defparam ram_block1a63.port_b_first_address = 0;
defparam ram_block1a63.port_b_first_bit_number = 63;
defparam ram_block1a63.port_b_last_address = 8191;
defparam ram_block1a63.port_b_logical_ram_depth = 16384;
defparam ram_block1a63.port_b_logical_ram_width = 64;
defparam ram_block1a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a63.port_b_read_enable_clock = "clock1";
defparam ram_block1a63.port_b_write_enable_clock = "clock1";
defparam ram_block1a63.ram_block_type = "auto";
defparam ram_block1a63.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a63.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a63.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block1a63.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

dffeas \address_reg_a[0] (
	.clk(clock1),
	.d(address_a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken0),
	.q(\address_reg_a[0]~q ),
	.prn(vcc));
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";

dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(address_b[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clocken1),
	.q(\address_reg_b[0]~q ),
	.prn(vcc));
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";

endmodule

module qtestpd_decode_d0b (
	eq_node_1,
	eq_node_0,
	onchip_memory2_0_s1_address_13,
	onchip_memory2_0_s1_chipselect,
	onchip_memory2_0_s1_write)/* synthesis synthesis_greybox=0 */;
output 	eq_node_1;
output 	eq_node_0;
input 	onchip_memory2_0_s1_address_13;
input 	onchip_memory2_0_s1_chipselect;
input 	onchip_memory2_0_s1_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneiv_lcell_comb \eq_node[1]~0 (
	.dataa(onchip_memory2_0_s1_address_13),
	.datab(onchip_memory2_0_s1_chipselect),
	.datac(onchip_memory2_0_s1_write),
	.datad(gnd),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
defparam \eq_node[1]~0 .lut_mask = 16'h8080;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \eq_node[0]~1 (
	.dataa(onchip_memory2_0_s1_chipselect),
	.datab(onchip_memory2_0_s1_write),
	.datac(gnd),
	.datad(onchip_memory2_0_s1_address_13),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
defparam \eq_node[0]~1 .lut_mask = 16'h0088;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";

endmodule

module qtestpd_decode_d0b_1 (
	eq_node_1,
	eq_node_0,
	onchip_memory2_0_s2_address_13,
	onchip_memory2_0_s2_chipselect,
	onchip_memory2_0_s2_write)/* synthesis synthesis_greybox=0 */;
output 	eq_node_1;
output 	eq_node_0;
input 	onchip_memory2_0_s2_address_13;
input 	onchip_memory2_0_s2_chipselect;
input 	onchip_memory2_0_s2_write;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneiv_lcell_comb \eq_node[1]~0 (
	.dataa(onchip_memory2_0_s2_address_13),
	.datab(onchip_memory2_0_s2_chipselect),
	.datac(onchip_memory2_0_s2_write),
	.datad(gnd),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
defparam \eq_node[1]~0 .lut_mask = 16'h8080;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \eq_node[0]~1 (
	.dataa(onchip_memory2_0_s2_chipselect),
	.datab(onchip_memory2_0_s2_write),
	.datac(gnd),
	.datad(onchip_memory2_0_s2_address_13),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
defparam \eq_node[0]~1 .lut_mask = 16'h0088;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";

endmodule

module qtestpd_mux_fsb (
	ram_block1a64,
	ram_block1a0,
	ram_block1a65,
	ram_block1a1,
	ram_block1a66,
	ram_block1a2,
	ram_block1a67,
	ram_block1a3,
	ram_block1a68,
	ram_block1a4,
	ram_block1a69,
	ram_block1a5,
	ram_block1a70,
	ram_block1a6,
	ram_block1a71,
	ram_block1a7,
	ram_block1a72,
	ram_block1a8,
	ram_block1a73,
	ram_block1a9,
	ram_block1a74,
	ram_block1a10,
	ram_block1a75,
	ram_block1a11,
	ram_block1a76,
	ram_block1a12,
	ram_block1a77,
	ram_block1a13,
	ram_block1a78,
	ram_block1a14,
	ram_block1a79,
	ram_block1a15,
	ram_block1a80,
	ram_block1a16,
	ram_block1a81,
	ram_block1a17,
	ram_block1a82,
	ram_block1a18,
	ram_block1a83,
	ram_block1a19,
	ram_block1a84,
	ram_block1a20,
	ram_block1a85,
	ram_block1a21,
	ram_block1a86,
	ram_block1a22,
	ram_block1a87,
	ram_block1a23,
	ram_block1a88,
	ram_block1a24,
	ram_block1a89,
	ram_block1a25,
	ram_block1a90,
	ram_block1a26,
	ram_block1a91,
	ram_block1a27,
	ram_block1a92,
	ram_block1a28,
	ram_block1a93,
	ram_block1a29,
	ram_block1a94,
	ram_block1a30,
	ram_block1a95,
	ram_block1a31,
	ram_block1a96,
	ram_block1a32,
	ram_block1a97,
	ram_block1a33,
	ram_block1a98,
	ram_block1a34,
	ram_block1a99,
	ram_block1a35,
	ram_block1a100,
	ram_block1a36,
	ram_block1a101,
	ram_block1a37,
	ram_block1a102,
	ram_block1a38,
	ram_block1a103,
	ram_block1a39,
	ram_block1a104,
	ram_block1a40,
	ram_block1a105,
	ram_block1a41,
	ram_block1a106,
	ram_block1a42,
	ram_block1a107,
	ram_block1a43,
	ram_block1a108,
	ram_block1a44,
	ram_block1a109,
	ram_block1a45,
	ram_block1a110,
	ram_block1a46,
	ram_block1a111,
	ram_block1a47,
	ram_block1a112,
	ram_block1a48,
	ram_block1a113,
	ram_block1a49,
	ram_block1a114,
	ram_block1a50,
	ram_block1a115,
	ram_block1a51,
	ram_block1a116,
	ram_block1a52,
	ram_block1a117,
	ram_block1a53,
	ram_block1a118,
	ram_block1a54,
	ram_block1a119,
	ram_block1a55,
	ram_block1a120,
	ram_block1a56,
	ram_block1a121,
	ram_block1a57,
	ram_block1a122,
	ram_block1a58,
	ram_block1a123,
	ram_block1a59,
	ram_block1a124,
	ram_block1a60,
	ram_block1a125,
	ram_block1a61,
	ram_block1a126,
	ram_block1a62,
	ram_block1a127,
	ram_block1a63,
	address_reg_a_0,
	result_node_0,
	result_node_1,
	result_node_2,
	result_node_3,
	result_node_4,
	result_node_5,
	result_node_6,
	result_node_7,
	result_node_8,
	result_node_9,
	result_node_10,
	result_node_11,
	result_node_12,
	result_node_13,
	result_node_14,
	result_node_15,
	result_node_16,
	result_node_17,
	result_node_18,
	result_node_19,
	result_node_20,
	result_node_21,
	result_node_22,
	result_node_23,
	result_node_24,
	result_node_25,
	result_node_26,
	result_node_27,
	result_node_28,
	result_node_29,
	result_node_30,
	result_node_31,
	result_node_32,
	result_node_33,
	result_node_34,
	result_node_35,
	result_node_36,
	result_node_37,
	result_node_38,
	result_node_39,
	result_node_40,
	result_node_41,
	result_node_42,
	result_node_43,
	result_node_44,
	result_node_45,
	result_node_46,
	result_node_47,
	result_node_48,
	result_node_49,
	result_node_50,
	result_node_51,
	result_node_52,
	result_node_53,
	result_node_54,
	result_node_55,
	result_node_56,
	result_node_57,
	result_node_58,
	result_node_59,
	result_node_60,
	result_node_61,
	result_node_62,
	result_node_63)/* synthesis synthesis_greybox=0 */;
input 	ram_block1a64;
input 	ram_block1a0;
input 	ram_block1a65;
input 	ram_block1a1;
input 	ram_block1a66;
input 	ram_block1a2;
input 	ram_block1a67;
input 	ram_block1a3;
input 	ram_block1a68;
input 	ram_block1a4;
input 	ram_block1a69;
input 	ram_block1a5;
input 	ram_block1a70;
input 	ram_block1a6;
input 	ram_block1a71;
input 	ram_block1a7;
input 	ram_block1a72;
input 	ram_block1a8;
input 	ram_block1a73;
input 	ram_block1a9;
input 	ram_block1a74;
input 	ram_block1a10;
input 	ram_block1a75;
input 	ram_block1a11;
input 	ram_block1a76;
input 	ram_block1a12;
input 	ram_block1a77;
input 	ram_block1a13;
input 	ram_block1a78;
input 	ram_block1a14;
input 	ram_block1a79;
input 	ram_block1a15;
input 	ram_block1a80;
input 	ram_block1a16;
input 	ram_block1a81;
input 	ram_block1a17;
input 	ram_block1a82;
input 	ram_block1a18;
input 	ram_block1a83;
input 	ram_block1a19;
input 	ram_block1a84;
input 	ram_block1a20;
input 	ram_block1a85;
input 	ram_block1a21;
input 	ram_block1a86;
input 	ram_block1a22;
input 	ram_block1a87;
input 	ram_block1a23;
input 	ram_block1a88;
input 	ram_block1a24;
input 	ram_block1a89;
input 	ram_block1a25;
input 	ram_block1a90;
input 	ram_block1a26;
input 	ram_block1a91;
input 	ram_block1a27;
input 	ram_block1a92;
input 	ram_block1a28;
input 	ram_block1a93;
input 	ram_block1a29;
input 	ram_block1a94;
input 	ram_block1a30;
input 	ram_block1a95;
input 	ram_block1a31;
input 	ram_block1a96;
input 	ram_block1a32;
input 	ram_block1a97;
input 	ram_block1a33;
input 	ram_block1a98;
input 	ram_block1a34;
input 	ram_block1a99;
input 	ram_block1a35;
input 	ram_block1a100;
input 	ram_block1a36;
input 	ram_block1a101;
input 	ram_block1a37;
input 	ram_block1a102;
input 	ram_block1a38;
input 	ram_block1a103;
input 	ram_block1a39;
input 	ram_block1a104;
input 	ram_block1a40;
input 	ram_block1a105;
input 	ram_block1a41;
input 	ram_block1a106;
input 	ram_block1a42;
input 	ram_block1a107;
input 	ram_block1a43;
input 	ram_block1a108;
input 	ram_block1a44;
input 	ram_block1a109;
input 	ram_block1a45;
input 	ram_block1a110;
input 	ram_block1a46;
input 	ram_block1a111;
input 	ram_block1a47;
input 	ram_block1a112;
input 	ram_block1a48;
input 	ram_block1a113;
input 	ram_block1a49;
input 	ram_block1a114;
input 	ram_block1a50;
input 	ram_block1a115;
input 	ram_block1a51;
input 	ram_block1a116;
input 	ram_block1a52;
input 	ram_block1a117;
input 	ram_block1a53;
input 	ram_block1a118;
input 	ram_block1a54;
input 	ram_block1a119;
input 	ram_block1a55;
input 	ram_block1a120;
input 	ram_block1a56;
input 	ram_block1a121;
input 	ram_block1a57;
input 	ram_block1a122;
input 	ram_block1a58;
input 	ram_block1a123;
input 	ram_block1a59;
input 	ram_block1a124;
input 	ram_block1a60;
input 	ram_block1a125;
input 	ram_block1a61;
input 	ram_block1a126;
input 	ram_block1a62;
input 	ram_block1a127;
input 	ram_block1a63;
input 	address_reg_a_0;
output 	result_node_0;
output 	result_node_1;
output 	result_node_2;
output 	result_node_3;
output 	result_node_4;
output 	result_node_5;
output 	result_node_6;
output 	result_node_7;
output 	result_node_8;
output 	result_node_9;
output 	result_node_10;
output 	result_node_11;
output 	result_node_12;
output 	result_node_13;
output 	result_node_14;
output 	result_node_15;
output 	result_node_16;
output 	result_node_17;
output 	result_node_18;
output 	result_node_19;
output 	result_node_20;
output 	result_node_21;
output 	result_node_22;
output 	result_node_23;
output 	result_node_24;
output 	result_node_25;
output 	result_node_26;
output 	result_node_27;
output 	result_node_28;
output 	result_node_29;
output 	result_node_30;
output 	result_node_31;
output 	result_node_32;
output 	result_node_33;
output 	result_node_34;
output 	result_node_35;
output 	result_node_36;
output 	result_node_37;
output 	result_node_38;
output 	result_node_39;
output 	result_node_40;
output 	result_node_41;
output 	result_node_42;
output 	result_node_43;
output 	result_node_44;
output 	result_node_45;
output 	result_node_46;
output 	result_node_47;
output 	result_node_48;
output 	result_node_49;
output 	result_node_50;
output 	result_node_51;
output 	result_node_52;
output 	result_node_53;
output 	result_node_54;
output 	result_node_55;
output 	result_node_56;
output 	result_node_57;
output 	result_node_58;
output 	result_node_59;
output 	result_node_60;
output 	result_node_61;
output 	result_node_62;
output 	result_node_63;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneiv_lcell_comb \result_node[0]~0 (
	.dataa(ram_block1a64),
	.datab(ram_block1a0),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_0),
	.cout());
defparam \result_node[0]~0 .lut_mask = 16'hAACC;
defparam \result_node[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[1]~1 (
	.dataa(ram_block1a65),
	.datab(ram_block1a1),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_1),
	.cout());
defparam \result_node[1]~1 .lut_mask = 16'hAACC;
defparam \result_node[1]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[2]~2 (
	.dataa(ram_block1a66),
	.datab(ram_block1a2),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_2),
	.cout());
defparam \result_node[2]~2 .lut_mask = 16'hAACC;
defparam \result_node[2]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[3]~3 (
	.dataa(ram_block1a67),
	.datab(ram_block1a3),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_3),
	.cout());
defparam \result_node[3]~3 .lut_mask = 16'hAACC;
defparam \result_node[3]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[4]~4 (
	.dataa(ram_block1a68),
	.datab(ram_block1a4),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_4),
	.cout());
defparam \result_node[4]~4 .lut_mask = 16'hAACC;
defparam \result_node[4]~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[5]~5 (
	.dataa(ram_block1a69),
	.datab(ram_block1a5),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_5),
	.cout());
defparam \result_node[5]~5 .lut_mask = 16'hAACC;
defparam \result_node[5]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[6]~6 (
	.dataa(ram_block1a70),
	.datab(ram_block1a6),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_6),
	.cout());
defparam \result_node[6]~6 .lut_mask = 16'hAACC;
defparam \result_node[6]~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[7]~7 (
	.dataa(ram_block1a71),
	.datab(ram_block1a7),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_7),
	.cout());
defparam \result_node[7]~7 .lut_mask = 16'hAACC;
defparam \result_node[7]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[8]~8 (
	.dataa(ram_block1a72),
	.datab(ram_block1a8),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_8),
	.cout());
defparam \result_node[8]~8 .lut_mask = 16'hAACC;
defparam \result_node[8]~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[9]~9 (
	.dataa(ram_block1a73),
	.datab(ram_block1a9),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_9),
	.cout());
defparam \result_node[9]~9 .lut_mask = 16'hAACC;
defparam \result_node[9]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[10]~10 (
	.dataa(ram_block1a74),
	.datab(ram_block1a10),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_10),
	.cout());
defparam \result_node[10]~10 .lut_mask = 16'hAACC;
defparam \result_node[10]~10 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[11]~11 (
	.dataa(ram_block1a75),
	.datab(ram_block1a11),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_11),
	.cout());
defparam \result_node[11]~11 .lut_mask = 16'hAACC;
defparam \result_node[11]~11 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[12]~12 (
	.dataa(ram_block1a76),
	.datab(ram_block1a12),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_12),
	.cout());
defparam \result_node[12]~12 .lut_mask = 16'hAACC;
defparam \result_node[12]~12 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[13]~13 (
	.dataa(ram_block1a77),
	.datab(ram_block1a13),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_13),
	.cout());
defparam \result_node[13]~13 .lut_mask = 16'hAACC;
defparam \result_node[13]~13 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[14]~14 (
	.dataa(ram_block1a78),
	.datab(ram_block1a14),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_14),
	.cout());
defparam \result_node[14]~14 .lut_mask = 16'hAACC;
defparam \result_node[14]~14 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[15]~15 (
	.dataa(ram_block1a79),
	.datab(ram_block1a15),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_15),
	.cout());
defparam \result_node[15]~15 .lut_mask = 16'hAACC;
defparam \result_node[15]~15 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[16]~16 (
	.dataa(ram_block1a80),
	.datab(ram_block1a16),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_16),
	.cout());
defparam \result_node[16]~16 .lut_mask = 16'hAACC;
defparam \result_node[16]~16 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[17]~17 (
	.dataa(ram_block1a81),
	.datab(ram_block1a17),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_17),
	.cout());
defparam \result_node[17]~17 .lut_mask = 16'hAACC;
defparam \result_node[17]~17 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[18]~18 (
	.dataa(ram_block1a82),
	.datab(ram_block1a18),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_18),
	.cout());
defparam \result_node[18]~18 .lut_mask = 16'hAACC;
defparam \result_node[18]~18 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[19]~19 (
	.dataa(ram_block1a83),
	.datab(ram_block1a19),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_19),
	.cout());
defparam \result_node[19]~19 .lut_mask = 16'hAACC;
defparam \result_node[19]~19 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[20]~20 (
	.dataa(ram_block1a84),
	.datab(ram_block1a20),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_20),
	.cout());
defparam \result_node[20]~20 .lut_mask = 16'hAACC;
defparam \result_node[20]~20 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[21]~21 (
	.dataa(ram_block1a85),
	.datab(ram_block1a21),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_21),
	.cout());
defparam \result_node[21]~21 .lut_mask = 16'hAACC;
defparam \result_node[21]~21 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[22]~22 (
	.dataa(ram_block1a86),
	.datab(ram_block1a22),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_22),
	.cout());
defparam \result_node[22]~22 .lut_mask = 16'hAACC;
defparam \result_node[22]~22 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[23]~23 (
	.dataa(ram_block1a87),
	.datab(ram_block1a23),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_23),
	.cout());
defparam \result_node[23]~23 .lut_mask = 16'hAACC;
defparam \result_node[23]~23 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[24]~24 (
	.dataa(ram_block1a88),
	.datab(ram_block1a24),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_24),
	.cout());
defparam \result_node[24]~24 .lut_mask = 16'hAACC;
defparam \result_node[24]~24 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[25]~25 (
	.dataa(ram_block1a89),
	.datab(ram_block1a25),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_25),
	.cout());
defparam \result_node[25]~25 .lut_mask = 16'hAACC;
defparam \result_node[25]~25 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[26]~26 (
	.dataa(ram_block1a90),
	.datab(ram_block1a26),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_26),
	.cout());
defparam \result_node[26]~26 .lut_mask = 16'hAACC;
defparam \result_node[26]~26 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[27]~27 (
	.dataa(ram_block1a91),
	.datab(ram_block1a27),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_27),
	.cout());
defparam \result_node[27]~27 .lut_mask = 16'hAACC;
defparam \result_node[27]~27 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[28]~28 (
	.dataa(ram_block1a92),
	.datab(ram_block1a28),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_28),
	.cout());
defparam \result_node[28]~28 .lut_mask = 16'hAACC;
defparam \result_node[28]~28 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[29]~29 (
	.dataa(ram_block1a93),
	.datab(ram_block1a29),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_29),
	.cout());
defparam \result_node[29]~29 .lut_mask = 16'hAACC;
defparam \result_node[29]~29 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[30]~30 (
	.dataa(ram_block1a94),
	.datab(ram_block1a30),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_30),
	.cout());
defparam \result_node[30]~30 .lut_mask = 16'hAACC;
defparam \result_node[30]~30 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[31]~31 (
	.dataa(ram_block1a95),
	.datab(ram_block1a31),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_31),
	.cout());
defparam \result_node[31]~31 .lut_mask = 16'hAACC;
defparam \result_node[31]~31 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[32]~32 (
	.dataa(ram_block1a96),
	.datab(ram_block1a32),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_32),
	.cout());
defparam \result_node[32]~32 .lut_mask = 16'hAACC;
defparam \result_node[32]~32 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[33]~33 (
	.dataa(ram_block1a97),
	.datab(ram_block1a33),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_33),
	.cout());
defparam \result_node[33]~33 .lut_mask = 16'hAACC;
defparam \result_node[33]~33 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[34]~34 (
	.dataa(ram_block1a98),
	.datab(ram_block1a34),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_34),
	.cout());
defparam \result_node[34]~34 .lut_mask = 16'hAACC;
defparam \result_node[34]~34 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[35]~35 (
	.dataa(ram_block1a99),
	.datab(ram_block1a35),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_35),
	.cout());
defparam \result_node[35]~35 .lut_mask = 16'hAACC;
defparam \result_node[35]~35 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[36]~36 (
	.dataa(ram_block1a100),
	.datab(ram_block1a36),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_36),
	.cout());
defparam \result_node[36]~36 .lut_mask = 16'hAACC;
defparam \result_node[36]~36 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[37]~37 (
	.dataa(ram_block1a101),
	.datab(ram_block1a37),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_37),
	.cout());
defparam \result_node[37]~37 .lut_mask = 16'hAACC;
defparam \result_node[37]~37 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[38]~38 (
	.dataa(ram_block1a102),
	.datab(ram_block1a38),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_38),
	.cout());
defparam \result_node[38]~38 .lut_mask = 16'hAACC;
defparam \result_node[38]~38 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[39]~39 (
	.dataa(ram_block1a103),
	.datab(ram_block1a39),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_39),
	.cout());
defparam \result_node[39]~39 .lut_mask = 16'hAACC;
defparam \result_node[39]~39 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[40]~40 (
	.dataa(ram_block1a104),
	.datab(ram_block1a40),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_40),
	.cout());
defparam \result_node[40]~40 .lut_mask = 16'hAACC;
defparam \result_node[40]~40 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[41]~41 (
	.dataa(ram_block1a105),
	.datab(ram_block1a41),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_41),
	.cout());
defparam \result_node[41]~41 .lut_mask = 16'hAACC;
defparam \result_node[41]~41 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[42]~42 (
	.dataa(ram_block1a106),
	.datab(ram_block1a42),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_42),
	.cout());
defparam \result_node[42]~42 .lut_mask = 16'hAACC;
defparam \result_node[42]~42 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[43]~43 (
	.dataa(ram_block1a107),
	.datab(ram_block1a43),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_43),
	.cout());
defparam \result_node[43]~43 .lut_mask = 16'hAACC;
defparam \result_node[43]~43 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[44]~44 (
	.dataa(ram_block1a108),
	.datab(ram_block1a44),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_44),
	.cout());
defparam \result_node[44]~44 .lut_mask = 16'hAACC;
defparam \result_node[44]~44 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[45]~45 (
	.dataa(ram_block1a109),
	.datab(ram_block1a45),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_45),
	.cout());
defparam \result_node[45]~45 .lut_mask = 16'hAACC;
defparam \result_node[45]~45 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[46]~46 (
	.dataa(ram_block1a110),
	.datab(ram_block1a46),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_46),
	.cout());
defparam \result_node[46]~46 .lut_mask = 16'hAACC;
defparam \result_node[46]~46 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[47]~47 (
	.dataa(ram_block1a111),
	.datab(ram_block1a47),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_47),
	.cout());
defparam \result_node[47]~47 .lut_mask = 16'hAACC;
defparam \result_node[47]~47 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[48]~48 (
	.dataa(ram_block1a112),
	.datab(ram_block1a48),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_48),
	.cout());
defparam \result_node[48]~48 .lut_mask = 16'hAACC;
defparam \result_node[48]~48 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[49]~49 (
	.dataa(ram_block1a113),
	.datab(ram_block1a49),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_49),
	.cout());
defparam \result_node[49]~49 .lut_mask = 16'hAACC;
defparam \result_node[49]~49 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[50]~50 (
	.dataa(ram_block1a114),
	.datab(ram_block1a50),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_50),
	.cout());
defparam \result_node[50]~50 .lut_mask = 16'hAACC;
defparam \result_node[50]~50 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[51]~51 (
	.dataa(ram_block1a115),
	.datab(ram_block1a51),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_51),
	.cout());
defparam \result_node[51]~51 .lut_mask = 16'hAACC;
defparam \result_node[51]~51 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[52]~52 (
	.dataa(ram_block1a116),
	.datab(ram_block1a52),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_52),
	.cout());
defparam \result_node[52]~52 .lut_mask = 16'hAACC;
defparam \result_node[52]~52 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[53]~53 (
	.dataa(ram_block1a117),
	.datab(ram_block1a53),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_53),
	.cout());
defparam \result_node[53]~53 .lut_mask = 16'hAACC;
defparam \result_node[53]~53 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[54]~54 (
	.dataa(ram_block1a118),
	.datab(ram_block1a54),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_54),
	.cout());
defparam \result_node[54]~54 .lut_mask = 16'hAACC;
defparam \result_node[54]~54 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[55]~55 (
	.dataa(ram_block1a119),
	.datab(ram_block1a55),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_55),
	.cout());
defparam \result_node[55]~55 .lut_mask = 16'hAACC;
defparam \result_node[55]~55 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[56]~56 (
	.dataa(ram_block1a120),
	.datab(ram_block1a56),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_56),
	.cout());
defparam \result_node[56]~56 .lut_mask = 16'hAACC;
defparam \result_node[56]~56 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[57]~57 (
	.dataa(ram_block1a121),
	.datab(ram_block1a57),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_57),
	.cout());
defparam \result_node[57]~57 .lut_mask = 16'hAACC;
defparam \result_node[57]~57 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[58]~58 (
	.dataa(ram_block1a122),
	.datab(ram_block1a58),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_58),
	.cout());
defparam \result_node[58]~58 .lut_mask = 16'hAACC;
defparam \result_node[58]~58 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[59]~59 (
	.dataa(ram_block1a123),
	.datab(ram_block1a59),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_59),
	.cout());
defparam \result_node[59]~59 .lut_mask = 16'hAACC;
defparam \result_node[59]~59 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[60]~60 (
	.dataa(ram_block1a124),
	.datab(ram_block1a60),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_60),
	.cout());
defparam \result_node[60]~60 .lut_mask = 16'hAACC;
defparam \result_node[60]~60 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[61]~61 (
	.dataa(ram_block1a125),
	.datab(ram_block1a61),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_61),
	.cout());
defparam \result_node[61]~61 .lut_mask = 16'hAACC;
defparam \result_node[61]~61 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[62]~62 (
	.dataa(ram_block1a126),
	.datab(ram_block1a62),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_62),
	.cout());
defparam \result_node[62]~62 .lut_mask = 16'hAACC;
defparam \result_node[62]~62 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[63]~63 (
	.dataa(ram_block1a127),
	.datab(ram_block1a63),
	.datac(gnd),
	.datad(address_reg_a_0),
	.cin(gnd),
	.combout(result_node_63),
	.cout());
defparam \result_node[63]~63 .lut_mask = 16'hAACC;
defparam \result_node[63]~63 .sum_lutc_input = "datac";

endmodule

module qtestpd_mux_fsb_1 (
	ram_block1a64,
	ram_block1a0,
	ram_block1a65,
	ram_block1a1,
	ram_block1a66,
	ram_block1a2,
	ram_block1a67,
	ram_block1a3,
	ram_block1a68,
	ram_block1a4,
	ram_block1a69,
	ram_block1a5,
	ram_block1a70,
	ram_block1a6,
	ram_block1a71,
	ram_block1a7,
	ram_block1a72,
	ram_block1a8,
	ram_block1a73,
	ram_block1a9,
	ram_block1a74,
	ram_block1a10,
	ram_block1a75,
	ram_block1a11,
	ram_block1a76,
	ram_block1a12,
	ram_block1a77,
	ram_block1a13,
	ram_block1a78,
	ram_block1a14,
	ram_block1a79,
	ram_block1a15,
	ram_block1a80,
	ram_block1a16,
	ram_block1a81,
	ram_block1a17,
	ram_block1a82,
	ram_block1a18,
	ram_block1a83,
	ram_block1a19,
	ram_block1a84,
	ram_block1a20,
	ram_block1a85,
	ram_block1a21,
	ram_block1a86,
	ram_block1a22,
	ram_block1a87,
	ram_block1a23,
	ram_block1a88,
	ram_block1a24,
	ram_block1a89,
	ram_block1a25,
	ram_block1a90,
	ram_block1a26,
	ram_block1a91,
	ram_block1a27,
	ram_block1a92,
	ram_block1a28,
	ram_block1a93,
	ram_block1a29,
	ram_block1a94,
	ram_block1a30,
	ram_block1a95,
	ram_block1a31,
	ram_block1a96,
	ram_block1a32,
	ram_block1a97,
	ram_block1a33,
	ram_block1a98,
	ram_block1a34,
	ram_block1a99,
	ram_block1a35,
	ram_block1a100,
	ram_block1a36,
	ram_block1a101,
	ram_block1a37,
	ram_block1a102,
	ram_block1a38,
	ram_block1a103,
	ram_block1a39,
	ram_block1a104,
	ram_block1a40,
	ram_block1a105,
	ram_block1a41,
	ram_block1a106,
	ram_block1a42,
	ram_block1a107,
	ram_block1a43,
	ram_block1a108,
	ram_block1a44,
	ram_block1a109,
	ram_block1a45,
	ram_block1a110,
	ram_block1a46,
	ram_block1a111,
	ram_block1a47,
	ram_block1a112,
	ram_block1a48,
	ram_block1a113,
	ram_block1a49,
	ram_block1a114,
	ram_block1a50,
	ram_block1a115,
	ram_block1a51,
	ram_block1a116,
	ram_block1a52,
	ram_block1a117,
	ram_block1a53,
	ram_block1a118,
	ram_block1a54,
	ram_block1a119,
	ram_block1a55,
	ram_block1a120,
	ram_block1a56,
	ram_block1a121,
	ram_block1a57,
	ram_block1a122,
	ram_block1a58,
	ram_block1a123,
	ram_block1a59,
	ram_block1a124,
	ram_block1a60,
	ram_block1a125,
	ram_block1a61,
	ram_block1a126,
	ram_block1a62,
	ram_block1a127,
	ram_block1a63,
	address_reg_b_0,
	result_node_0,
	result_node_1,
	result_node_2,
	result_node_3,
	result_node_4,
	result_node_5,
	result_node_6,
	result_node_7,
	result_node_8,
	result_node_9,
	result_node_10,
	result_node_11,
	result_node_12,
	result_node_13,
	result_node_14,
	result_node_15,
	result_node_16,
	result_node_17,
	result_node_18,
	result_node_19,
	result_node_20,
	result_node_21,
	result_node_22,
	result_node_23,
	result_node_24,
	result_node_25,
	result_node_26,
	result_node_27,
	result_node_28,
	result_node_29,
	result_node_30,
	result_node_31,
	result_node_32,
	result_node_33,
	result_node_34,
	result_node_35,
	result_node_36,
	result_node_37,
	result_node_38,
	result_node_39,
	result_node_40,
	result_node_41,
	result_node_42,
	result_node_43,
	result_node_44,
	result_node_45,
	result_node_46,
	result_node_47,
	result_node_48,
	result_node_49,
	result_node_50,
	result_node_51,
	result_node_52,
	result_node_53,
	result_node_54,
	result_node_55,
	result_node_56,
	result_node_57,
	result_node_58,
	result_node_59,
	result_node_60,
	result_node_61,
	result_node_62,
	result_node_63)/* synthesis synthesis_greybox=0 */;
input 	ram_block1a64;
input 	ram_block1a0;
input 	ram_block1a65;
input 	ram_block1a1;
input 	ram_block1a66;
input 	ram_block1a2;
input 	ram_block1a67;
input 	ram_block1a3;
input 	ram_block1a68;
input 	ram_block1a4;
input 	ram_block1a69;
input 	ram_block1a5;
input 	ram_block1a70;
input 	ram_block1a6;
input 	ram_block1a71;
input 	ram_block1a7;
input 	ram_block1a72;
input 	ram_block1a8;
input 	ram_block1a73;
input 	ram_block1a9;
input 	ram_block1a74;
input 	ram_block1a10;
input 	ram_block1a75;
input 	ram_block1a11;
input 	ram_block1a76;
input 	ram_block1a12;
input 	ram_block1a77;
input 	ram_block1a13;
input 	ram_block1a78;
input 	ram_block1a14;
input 	ram_block1a79;
input 	ram_block1a15;
input 	ram_block1a80;
input 	ram_block1a16;
input 	ram_block1a81;
input 	ram_block1a17;
input 	ram_block1a82;
input 	ram_block1a18;
input 	ram_block1a83;
input 	ram_block1a19;
input 	ram_block1a84;
input 	ram_block1a20;
input 	ram_block1a85;
input 	ram_block1a21;
input 	ram_block1a86;
input 	ram_block1a22;
input 	ram_block1a87;
input 	ram_block1a23;
input 	ram_block1a88;
input 	ram_block1a24;
input 	ram_block1a89;
input 	ram_block1a25;
input 	ram_block1a90;
input 	ram_block1a26;
input 	ram_block1a91;
input 	ram_block1a27;
input 	ram_block1a92;
input 	ram_block1a28;
input 	ram_block1a93;
input 	ram_block1a29;
input 	ram_block1a94;
input 	ram_block1a30;
input 	ram_block1a95;
input 	ram_block1a31;
input 	ram_block1a96;
input 	ram_block1a32;
input 	ram_block1a97;
input 	ram_block1a33;
input 	ram_block1a98;
input 	ram_block1a34;
input 	ram_block1a99;
input 	ram_block1a35;
input 	ram_block1a100;
input 	ram_block1a36;
input 	ram_block1a101;
input 	ram_block1a37;
input 	ram_block1a102;
input 	ram_block1a38;
input 	ram_block1a103;
input 	ram_block1a39;
input 	ram_block1a104;
input 	ram_block1a40;
input 	ram_block1a105;
input 	ram_block1a41;
input 	ram_block1a106;
input 	ram_block1a42;
input 	ram_block1a107;
input 	ram_block1a43;
input 	ram_block1a108;
input 	ram_block1a44;
input 	ram_block1a109;
input 	ram_block1a45;
input 	ram_block1a110;
input 	ram_block1a46;
input 	ram_block1a111;
input 	ram_block1a47;
input 	ram_block1a112;
input 	ram_block1a48;
input 	ram_block1a113;
input 	ram_block1a49;
input 	ram_block1a114;
input 	ram_block1a50;
input 	ram_block1a115;
input 	ram_block1a51;
input 	ram_block1a116;
input 	ram_block1a52;
input 	ram_block1a117;
input 	ram_block1a53;
input 	ram_block1a118;
input 	ram_block1a54;
input 	ram_block1a119;
input 	ram_block1a55;
input 	ram_block1a120;
input 	ram_block1a56;
input 	ram_block1a121;
input 	ram_block1a57;
input 	ram_block1a122;
input 	ram_block1a58;
input 	ram_block1a123;
input 	ram_block1a59;
input 	ram_block1a124;
input 	ram_block1a60;
input 	ram_block1a125;
input 	ram_block1a61;
input 	ram_block1a126;
input 	ram_block1a62;
input 	ram_block1a127;
input 	ram_block1a63;
input 	address_reg_b_0;
output 	result_node_0;
output 	result_node_1;
output 	result_node_2;
output 	result_node_3;
output 	result_node_4;
output 	result_node_5;
output 	result_node_6;
output 	result_node_7;
output 	result_node_8;
output 	result_node_9;
output 	result_node_10;
output 	result_node_11;
output 	result_node_12;
output 	result_node_13;
output 	result_node_14;
output 	result_node_15;
output 	result_node_16;
output 	result_node_17;
output 	result_node_18;
output 	result_node_19;
output 	result_node_20;
output 	result_node_21;
output 	result_node_22;
output 	result_node_23;
output 	result_node_24;
output 	result_node_25;
output 	result_node_26;
output 	result_node_27;
output 	result_node_28;
output 	result_node_29;
output 	result_node_30;
output 	result_node_31;
output 	result_node_32;
output 	result_node_33;
output 	result_node_34;
output 	result_node_35;
output 	result_node_36;
output 	result_node_37;
output 	result_node_38;
output 	result_node_39;
output 	result_node_40;
output 	result_node_41;
output 	result_node_42;
output 	result_node_43;
output 	result_node_44;
output 	result_node_45;
output 	result_node_46;
output 	result_node_47;
output 	result_node_48;
output 	result_node_49;
output 	result_node_50;
output 	result_node_51;
output 	result_node_52;
output 	result_node_53;
output 	result_node_54;
output 	result_node_55;
output 	result_node_56;
output 	result_node_57;
output 	result_node_58;
output 	result_node_59;
output 	result_node_60;
output 	result_node_61;
output 	result_node_62;
output 	result_node_63;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneiv_lcell_comb \result_node[0]~0 (
	.dataa(ram_block1a64),
	.datab(ram_block1a0),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_0),
	.cout());
defparam \result_node[0]~0 .lut_mask = 16'hAACC;
defparam \result_node[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[1]~1 (
	.dataa(ram_block1a65),
	.datab(ram_block1a1),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_1),
	.cout());
defparam \result_node[1]~1 .lut_mask = 16'hAACC;
defparam \result_node[1]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[2]~2 (
	.dataa(ram_block1a66),
	.datab(ram_block1a2),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_2),
	.cout());
defparam \result_node[2]~2 .lut_mask = 16'hAACC;
defparam \result_node[2]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[3]~3 (
	.dataa(ram_block1a67),
	.datab(ram_block1a3),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_3),
	.cout());
defparam \result_node[3]~3 .lut_mask = 16'hAACC;
defparam \result_node[3]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[4]~4 (
	.dataa(ram_block1a68),
	.datab(ram_block1a4),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_4),
	.cout());
defparam \result_node[4]~4 .lut_mask = 16'hAACC;
defparam \result_node[4]~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[5]~5 (
	.dataa(ram_block1a69),
	.datab(ram_block1a5),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_5),
	.cout());
defparam \result_node[5]~5 .lut_mask = 16'hAACC;
defparam \result_node[5]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[6]~6 (
	.dataa(ram_block1a70),
	.datab(ram_block1a6),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_6),
	.cout());
defparam \result_node[6]~6 .lut_mask = 16'hAACC;
defparam \result_node[6]~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[7]~7 (
	.dataa(ram_block1a71),
	.datab(ram_block1a7),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_7),
	.cout());
defparam \result_node[7]~7 .lut_mask = 16'hAACC;
defparam \result_node[7]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[8]~8 (
	.dataa(ram_block1a72),
	.datab(ram_block1a8),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_8),
	.cout());
defparam \result_node[8]~8 .lut_mask = 16'hAACC;
defparam \result_node[8]~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[9]~9 (
	.dataa(ram_block1a73),
	.datab(ram_block1a9),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_9),
	.cout());
defparam \result_node[9]~9 .lut_mask = 16'hAACC;
defparam \result_node[9]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[10]~10 (
	.dataa(ram_block1a74),
	.datab(ram_block1a10),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_10),
	.cout());
defparam \result_node[10]~10 .lut_mask = 16'hAACC;
defparam \result_node[10]~10 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[11]~11 (
	.dataa(ram_block1a75),
	.datab(ram_block1a11),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_11),
	.cout());
defparam \result_node[11]~11 .lut_mask = 16'hAACC;
defparam \result_node[11]~11 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[12]~12 (
	.dataa(ram_block1a76),
	.datab(ram_block1a12),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_12),
	.cout());
defparam \result_node[12]~12 .lut_mask = 16'hAACC;
defparam \result_node[12]~12 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[13]~13 (
	.dataa(ram_block1a77),
	.datab(ram_block1a13),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_13),
	.cout());
defparam \result_node[13]~13 .lut_mask = 16'hAACC;
defparam \result_node[13]~13 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[14]~14 (
	.dataa(ram_block1a78),
	.datab(ram_block1a14),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_14),
	.cout());
defparam \result_node[14]~14 .lut_mask = 16'hAACC;
defparam \result_node[14]~14 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[15]~15 (
	.dataa(ram_block1a79),
	.datab(ram_block1a15),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_15),
	.cout());
defparam \result_node[15]~15 .lut_mask = 16'hAACC;
defparam \result_node[15]~15 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[16]~16 (
	.dataa(ram_block1a80),
	.datab(ram_block1a16),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_16),
	.cout());
defparam \result_node[16]~16 .lut_mask = 16'hAACC;
defparam \result_node[16]~16 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[17]~17 (
	.dataa(ram_block1a81),
	.datab(ram_block1a17),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_17),
	.cout());
defparam \result_node[17]~17 .lut_mask = 16'hAACC;
defparam \result_node[17]~17 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[18]~18 (
	.dataa(ram_block1a82),
	.datab(ram_block1a18),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_18),
	.cout());
defparam \result_node[18]~18 .lut_mask = 16'hAACC;
defparam \result_node[18]~18 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[19]~19 (
	.dataa(ram_block1a83),
	.datab(ram_block1a19),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_19),
	.cout());
defparam \result_node[19]~19 .lut_mask = 16'hAACC;
defparam \result_node[19]~19 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[20]~20 (
	.dataa(ram_block1a84),
	.datab(ram_block1a20),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_20),
	.cout());
defparam \result_node[20]~20 .lut_mask = 16'hAACC;
defparam \result_node[20]~20 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[21]~21 (
	.dataa(ram_block1a85),
	.datab(ram_block1a21),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_21),
	.cout());
defparam \result_node[21]~21 .lut_mask = 16'hAACC;
defparam \result_node[21]~21 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[22]~22 (
	.dataa(ram_block1a86),
	.datab(ram_block1a22),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_22),
	.cout());
defparam \result_node[22]~22 .lut_mask = 16'hAACC;
defparam \result_node[22]~22 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[23]~23 (
	.dataa(ram_block1a87),
	.datab(ram_block1a23),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_23),
	.cout());
defparam \result_node[23]~23 .lut_mask = 16'hAACC;
defparam \result_node[23]~23 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[24]~24 (
	.dataa(ram_block1a88),
	.datab(ram_block1a24),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_24),
	.cout());
defparam \result_node[24]~24 .lut_mask = 16'hAACC;
defparam \result_node[24]~24 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[25]~25 (
	.dataa(ram_block1a89),
	.datab(ram_block1a25),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_25),
	.cout());
defparam \result_node[25]~25 .lut_mask = 16'hAACC;
defparam \result_node[25]~25 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[26]~26 (
	.dataa(ram_block1a90),
	.datab(ram_block1a26),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_26),
	.cout());
defparam \result_node[26]~26 .lut_mask = 16'hAACC;
defparam \result_node[26]~26 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[27]~27 (
	.dataa(ram_block1a91),
	.datab(ram_block1a27),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_27),
	.cout());
defparam \result_node[27]~27 .lut_mask = 16'hAACC;
defparam \result_node[27]~27 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[28]~28 (
	.dataa(ram_block1a92),
	.datab(ram_block1a28),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_28),
	.cout());
defparam \result_node[28]~28 .lut_mask = 16'hAACC;
defparam \result_node[28]~28 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[29]~29 (
	.dataa(ram_block1a93),
	.datab(ram_block1a29),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_29),
	.cout());
defparam \result_node[29]~29 .lut_mask = 16'hAACC;
defparam \result_node[29]~29 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[30]~30 (
	.dataa(ram_block1a94),
	.datab(ram_block1a30),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_30),
	.cout());
defparam \result_node[30]~30 .lut_mask = 16'hAACC;
defparam \result_node[30]~30 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[31]~31 (
	.dataa(ram_block1a95),
	.datab(ram_block1a31),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_31),
	.cout());
defparam \result_node[31]~31 .lut_mask = 16'hAACC;
defparam \result_node[31]~31 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[32]~32 (
	.dataa(ram_block1a96),
	.datab(ram_block1a32),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_32),
	.cout());
defparam \result_node[32]~32 .lut_mask = 16'hAACC;
defparam \result_node[32]~32 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[33]~33 (
	.dataa(ram_block1a97),
	.datab(ram_block1a33),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_33),
	.cout());
defparam \result_node[33]~33 .lut_mask = 16'hAACC;
defparam \result_node[33]~33 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[34]~34 (
	.dataa(ram_block1a98),
	.datab(ram_block1a34),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_34),
	.cout());
defparam \result_node[34]~34 .lut_mask = 16'hAACC;
defparam \result_node[34]~34 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[35]~35 (
	.dataa(ram_block1a99),
	.datab(ram_block1a35),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_35),
	.cout());
defparam \result_node[35]~35 .lut_mask = 16'hAACC;
defparam \result_node[35]~35 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[36]~36 (
	.dataa(ram_block1a100),
	.datab(ram_block1a36),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_36),
	.cout());
defparam \result_node[36]~36 .lut_mask = 16'hAACC;
defparam \result_node[36]~36 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[37]~37 (
	.dataa(ram_block1a101),
	.datab(ram_block1a37),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_37),
	.cout());
defparam \result_node[37]~37 .lut_mask = 16'hAACC;
defparam \result_node[37]~37 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[38]~38 (
	.dataa(ram_block1a102),
	.datab(ram_block1a38),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_38),
	.cout());
defparam \result_node[38]~38 .lut_mask = 16'hAACC;
defparam \result_node[38]~38 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[39]~39 (
	.dataa(ram_block1a103),
	.datab(ram_block1a39),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_39),
	.cout());
defparam \result_node[39]~39 .lut_mask = 16'hAACC;
defparam \result_node[39]~39 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[40]~40 (
	.dataa(ram_block1a104),
	.datab(ram_block1a40),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_40),
	.cout());
defparam \result_node[40]~40 .lut_mask = 16'hAACC;
defparam \result_node[40]~40 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[41]~41 (
	.dataa(ram_block1a105),
	.datab(ram_block1a41),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_41),
	.cout());
defparam \result_node[41]~41 .lut_mask = 16'hAACC;
defparam \result_node[41]~41 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[42]~42 (
	.dataa(ram_block1a106),
	.datab(ram_block1a42),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_42),
	.cout());
defparam \result_node[42]~42 .lut_mask = 16'hAACC;
defparam \result_node[42]~42 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[43]~43 (
	.dataa(ram_block1a107),
	.datab(ram_block1a43),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_43),
	.cout());
defparam \result_node[43]~43 .lut_mask = 16'hAACC;
defparam \result_node[43]~43 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[44]~44 (
	.dataa(ram_block1a108),
	.datab(ram_block1a44),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_44),
	.cout());
defparam \result_node[44]~44 .lut_mask = 16'hAACC;
defparam \result_node[44]~44 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[45]~45 (
	.dataa(ram_block1a109),
	.datab(ram_block1a45),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_45),
	.cout());
defparam \result_node[45]~45 .lut_mask = 16'hAACC;
defparam \result_node[45]~45 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[46]~46 (
	.dataa(ram_block1a110),
	.datab(ram_block1a46),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_46),
	.cout());
defparam \result_node[46]~46 .lut_mask = 16'hAACC;
defparam \result_node[46]~46 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[47]~47 (
	.dataa(ram_block1a111),
	.datab(ram_block1a47),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_47),
	.cout());
defparam \result_node[47]~47 .lut_mask = 16'hAACC;
defparam \result_node[47]~47 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[48]~48 (
	.dataa(ram_block1a112),
	.datab(ram_block1a48),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_48),
	.cout());
defparam \result_node[48]~48 .lut_mask = 16'hAACC;
defparam \result_node[48]~48 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[49]~49 (
	.dataa(ram_block1a113),
	.datab(ram_block1a49),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_49),
	.cout());
defparam \result_node[49]~49 .lut_mask = 16'hAACC;
defparam \result_node[49]~49 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[50]~50 (
	.dataa(ram_block1a114),
	.datab(ram_block1a50),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_50),
	.cout());
defparam \result_node[50]~50 .lut_mask = 16'hAACC;
defparam \result_node[50]~50 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[51]~51 (
	.dataa(ram_block1a115),
	.datab(ram_block1a51),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_51),
	.cout());
defparam \result_node[51]~51 .lut_mask = 16'hAACC;
defparam \result_node[51]~51 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[52]~52 (
	.dataa(ram_block1a116),
	.datab(ram_block1a52),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_52),
	.cout());
defparam \result_node[52]~52 .lut_mask = 16'hAACC;
defparam \result_node[52]~52 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[53]~53 (
	.dataa(ram_block1a117),
	.datab(ram_block1a53),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_53),
	.cout());
defparam \result_node[53]~53 .lut_mask = 16'hAACC;
defparam \result_node[53]~53 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[54]~54 (
	.dataa(ram_block1a118),
	.datab(ram_block1a54),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_54),
	.cout());
defparam \result_node[54]~54 .lut_mask = 16'hAACC;
defparam \result_node[54]~54 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[55]~55 (
	.dataa(ram_block1a119),
	.datab(ram_block1a55),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_55),
	.cout());
defparam \result_node[55]~55 .lut_mask = 16'hAACC;
defparam \result_node[55]~55 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[56]~56 (
	.dataa(ram_block1a120),
	.datab(ram_block1a56),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_56),
	.cout());
defparam \result_node[56]~56 .lut_mask = 16'hAACC;
defparam \result_node[56]~56 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[57]~57 (
	.dataa(ram_block1a121),
	.datab(ram_block1a57),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_57),
	.cout());
defparam \result_node[57]~57 .lut_mask = 16'hAACC;
defparam \result_node[57]~57 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[58]~58 (
	.dataa(ram_block1a122),
	.datab(ram_block1a58),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_58),
	.cout());
defparam \result_node[58]~58 .lut_mask = 16'hAACC;
defparam \result_node[58]~58 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[59]~59 (
	.dataa(ram_block1a123),
	.datab(ram_block1a59),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_59),
	.cout());
defparam \result_node[59]~59 .lut_mask = 16'hAACC;
defparam \result_node[59]~59 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[60]~60 (
	.dataa(ram_block1a124),
	.datab(ram_block1a60),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_60),
	.cout());
defparam \result_node[60]~60 .lut_mask = 16'hAACC;
defparam \result_node[60]~60 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[61]~61 (
	.dataa(ram_block1a125),
	.datab(ram_block1a61),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_61),
	.cout());
defparam \result_node[61]~61 .lut_mask = 16'hAACC;
defparam \result_node[61]~61 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[62]~62 (
	.dataa(ram_block1a126),
	.datab(ram_block1a62),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_62),
	.cout());
defparam \result_node[62]~62 .lut_mask = 16'hAACC;
defparam \result_node[62]~62 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \result_node[63]~63 (
	.dataa(ram_block1a127),
	.datab(ram_block1a63),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(result_node_63),
	.cout());
defparam \result_node[63]~63 .lut_mask = 16'hAACC;
defparam \result_node[63]~63 .sum_lutc_input = "datac";

endmodule
