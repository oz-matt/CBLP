// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"

// DATE "08/06/2019 23:31:21"

// 
// Device: Altera 5CSEBA6U23I7 Package UFBGA672
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module embedded_system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	ad9833_io_readdata,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
output 	[31:0] ad9833_io_readdata;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ad9833_comp_0|aif|fsync~q ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ;
wire \onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[2]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[10]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[18]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[26]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[7]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[23]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[15]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[31]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[29]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[13]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[28]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[12]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[27]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[11]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[25]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[9]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[24]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[8]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[6]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[14]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[22]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[30]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[5]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[21]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[4]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[20]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[3]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[19]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[1]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[17]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[0]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[16]~q ;
wire \ad9833_comp_0|aif|good_to_reset_go~q ;
wire \ad9833_comp_0|aif|send_complete~q ;
wire \ad9833_comp_0|aif|sclk~q ;
wire \ad9833_comp_0|aif|sdata~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[0]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[0]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[1]~q ;
wire \rst_controller|r_sync_rst~q ;
wire \mm_interconnect_0|ad9833_comp_0_avalon_slave_0_translator|wait_latency_counter[1]~q ;
wire \mm_interconnect_0|ad9833_comp_0_avalon_slave_0_translator|wait_latency_counter[0]~q ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_agent|hold_waitrequest~q ;
wire \nios2_qsys_0|d_address_offset_field[0]~q ;
wire \nios2_qsys_0|d_write~reg0_q ;
wire \nios2_qsys_0|d_address_tag_field[2]~q ;
wire \nios2_qsys_0|d_address_tag_field[1]~q ;
wire \nios2_qsys_0|d_address_tag_field[0]~q ;
wire \nios2_qsys_0|d_address_line_field[5]~q ;
wire \nios2_qsys_0|d_address_line_field[4]~q ;
wire \nios2_qsys_0|d_address_line_field[3]~q ;
wire \nios2_qsys_0|d_address_line_field[2]~q ;
wire \nios2_qsys_0|d_address_line_field[1]~q ;
wire \nios2_qsys_0|d_address_line_field[0]~q ;
wire \nios2_qsys_0|d_address_offset_field[2]~q ;
wire \nios2_qsys_0|d_address_offset_field[1]~q ;
wire \mm_interconnect_0|ad9833_comp_0_avalon_slave_0_agent|m0_write~0_combout ;
wire \nios2_qsys_0|d_writedata[11]~reg0_q ;
wire \nios2_qsys_0|d_byteenable[0]~reg0_q ;
wire \nios2_qsys_0|d_writedata[10]~reg0_q ;
wire \nios2_qsys_0|d_writedata[9]~reg0_q ;
wire \nios2_qsys_0|d_writedata[8]~reg0_q ;
wire \nios2_qsys_0|d_writedata[13]~reg0_q ;
wire \nios2_qsys_0|d_writedata[12]~reg0_q ;
wire \nios2_qsys_0|d_writedata[21]~reg0_q ;
wire \nios2_qsys_0|d_writedata[20]~reg0_q ;
wire \nios2_qsys_0|d_writedata[25]~reg0_q ;
wire \nios2_qsys_0|d_writedata[17]~reg0_q ;
wire \nios2_qsys_0|d_writedata[24]~reg0_q ;
wire \nios2_qsys_0|d_writedata[16]~reg0_q ;
wire \nios2_qsys_0|d_writedata[27]~reg0_q ;
wire \nios2_qsys_0|d_writedata[19]~reg0_q ;
wire \nios2_qsys_0|d_writedata[26]~reg0_q ;
wire \nios2_qsys_0|d_writedata[18]~reg0_q ;
wire \nios2_qsys_0|d_writedata[23]~reg0_q ;
wire \nios2_qsys_0|d_writedata[15]~reg0_q ;
wire \nios2_qsys_0|d_writedata[22]~reg0_q ;
wire \nios2_qsys_0|d_writedata[14]~reg0_q ;
wire \nios2_qsys_0|d_read~reg0_q ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_limiter|suppress_change_dest_id~0_combout ;
wire \mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_ocimem|waitrequest~q ;
wire \mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ;
wire \mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ;
wire \mm_interconnect_0|cmd_demux|WideOr0~combout ;
wire \mm_interconnect_0|nios2_qsys_0_data_master_agent|av_waitrequest~combout ;
wire \nios2_qsys_0|d_byteenable[1]~reg0_q ;
wire \nios2_qsys_0|d_writedata[2]~reg0_q ;
wire \nios2_qsys_0|d_writedata[0]~reg0_q ;
wire \nios2_qsys_0|d_writedata[3]~reg0_q ;
wire \nios2_qsys_0|d_writedata[1]~reg0_q ;
wire \nios2_qsys_0|hbreak_enabled~q ;
wire \nios2_qsys_0|i_read~reg0_q ;
wire \mm_interconnect_0|cmd_demux_001|src0_valid~0_combout ;
wire \nios2_qsys_0|ic_fill_tag[1]~q ;
wire \nios2_qsys_0|ic_fill_tag[0]~q ;
wire \nios2_qsys_0|ic_fill_line[6]~q ;
wire \mm_interconnect_0|router_001|Equal1~0_combout ;
wire \mm_interconnect_0|cmd_demux_001|src0_valid~1_combout ;
wire \mm_interconnect_0|cmd_demux|src1_valid~0_combout ;
wire \mm_interconnect_0|cmd_mux_001|saved_grant[1]~q ;
wire \mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent|rf_source_valid~0_combout ;
wire \mm_interconnect_0|cmd_demux_001|src1_valid~0_combout ;
wire \mm_interconnect_0|cmd_demux|src2_valid~2_combout ;
wire \mm_interconnect_0|cmd_mux_002|saved_grant[1]~q ;
wire \nios2_qsys_0|d_writedata[6]~reg0_q ;
wire \nios2_qsys_0|d_writedata[4]~reg0_q ;
wire \nios2_qsys_0|d_writedata[7]~reg0_q ;
wire \nios2_qsys_0|d_writedata[5]~reg0_q ;
wire \rst_controller|r_early_rst~q ;
wire \mm_interconnect_0|rsp_mux|WideOr1~combout ;
wire \mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|suppress_change_dest_id~0_combout ;
wire \mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ;
wire \mm_interconnect_0|cmd_demux_001|WideOr0~1_combout ;
wire \mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|nonposted_cmd_accepted~combout ;
wire \nios2_qsys_0|ic_fill_line[5]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~0_combout ;
wire \nios2_qsys_0|ic_fill_ap_offset[0]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[38]~combout ;
wire \nios2_qsys_0|ic_fill_line[1]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[42]~combout ;
wire \nios2_qsys_0|ic_fill_line[0]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[41]~combout ;
wire \nios2_qsys_0|ic_fill_ap_offset[2]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[40]~combout ;
wire \nios2_qsys_0|ic_fill_ap_offset[1]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[39]~combout ;
wire \nios2_qsys_0|ic_fill_line[4]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[45]~combout ;
wire \nios2_qsys_0|ic_fill_line[3]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[44]~combout ;
wire \nios2_qsys_0|ic_fill_line[2]~q ;
wire \mm_interconnect_0|cmd_mux_001|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[32]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~2_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~3_combout ;
wire \mm_interconnect_0|rsp_mux_001|WideOr1~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[2]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[10]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[18]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[26]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[7]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[23]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[15]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[31]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[29]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[13]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[28]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[12]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[27]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[11]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[25]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[9]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[24]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[8]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[6]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[14]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[22]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[30]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[5]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[21]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[4]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[20]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[3]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[19]~combout ;
wire \nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_oci_debug|resetrequest~q ;
wire \mm_interconnect_0|rsp_mux|src_data[1]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[17]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[0]~combout ;
wire \mm_interconnect_0|rsp_mux|src_data[16]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~4_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[5]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[3]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[1]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[4]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[2]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[28]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[31]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[27]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[29]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[30]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[0]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[23]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[26]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[22]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[24]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[25]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[16]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[15]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[13]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[14]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[12]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[11]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[8]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~0_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[38]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[39]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[40]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[41]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[42]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[43]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[44]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[45]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[46]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[47]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[32]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~1_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~2_combout ;
wire \nios2_qsys_0|d_byteenable[2]~reg0_q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~3_combout ;
wire \nios2_qsys_0|d_byteenable[3]~reg0_q ;
wire \mm_interconnect_0|cmd_mux_002|src_data[35]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[19]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~4_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~6_combout ;
wire \nios2_qsys_0|d_writedata[31]~reg0_q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~7_combout ;
wire \nios2_qsys_0|d_writedata[29]~reg0_q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~9_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[18]~combout ;
wire \nios2_qsys_0|d_writedata[28]~reg0_q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~11_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[17]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~20_combout ;
wire \nios2_qsys_0|d_writedata[30]~reg0_q ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~23_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[10]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~25_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[9]~combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_002|src_payload~31_combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[21]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[20]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[7]~combout ;
wire \mm_interconnect_0|rsp_mux_001|src_data[6]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~5_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[35]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~6_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~7_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[34]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~8_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~9_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~10_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~11_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~12_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~13_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~14_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~15_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~16_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~17_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~18_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~19_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~20_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~21_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_data[33]~combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~22_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~23_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~24_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~25_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~26_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~27_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~28_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~29_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~30_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~31_combout ;
wire \mm_interconnect_0|cmd_mux_001|src_payload~32_combout ;
wire \rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \clk_clk~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ;
wire \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|Equal2~2_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~q ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ;
wire \nabboc|pzdyqx_impl_inst|Equal2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ;
wire \nabboc|pzdyqx_impl_inst|comb~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ;
wire \nabboc|pzdyqx_impl_inst|sdr~combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ;
wire \nabboc|pzdyqx_impl_inst|dr_scan~combout ;
wire \nabboc|pzdyqx_impl_inst|KNOR6738~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \altera_internal_jtag~TDO ;


embedded_system_ad9833_avalon ad9833_comp_0(
	.fsync(\ad9833_comp_0|aif|fsync~q ),
	.good_to_reset_go(\ad9833_comp_0|aif|good_to_reset_go~q ),
	.send_complete(\ad9833_comp_0|aif|send_complete~q ),
	.sclk(\ad9833_comp_0|aif|sclk~q ),
	.sdata(\ad9833_comp_0|aif|sdata~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.wait_latency_counter_1(\mm_interconnect_0|ad9833_comp_0_avalon_slave_0_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|ad9833_comp_0_avalon_slave_0_translator|wait_latency_counter[0]~q ),
	.m0_write(\mm_interconnect_0|ad9833_comp_0_avalon_slave_0_agent|m0_write~0_combout ),
	.d_writedata_11(\nios2_qsys_0|d_writedata[11]~reg0_q ),
	.d_byteenable_0(\nios2_qsys_0|d_byteenable[0]~reg0_q ),
	.d_writedata_10(\nios2_qsys_0|d_writedata[10]~reg0_q ),
	.d_writedata_9(\nios2_qsys_0|d_writedata[9]~reg0_q ),
	.d_writedata_8(\nios2_qsys_0|d_writedata[8]~reg0_q ),
	.d_writedata_13(\nios2_qsys_0|d_writedata[13]~reg0_q ),
	.d_writedata_12(\nios2_qsys_0|d_writedata[12]~reg0_q ),
	.d_writedata_21(\nios2_qsys_0|d_writedata[21]~reg0_q ),
	.d_writedata_20(\nios2_qsys_0|d_writedata[20]~reg0_q ),
	.d_writedata_25(\nios2_qsys_0|d_writedata[25]~reg0_q ),
	.d_writedata_17(\nios2_qsys_0|d_writedata[17]~reg0_q ),
	.d_writedata_24(\nios2_qsys_0|d_writedata[24]~reg0_q ),
	.d_writedata_16(\nios2_qsys_0|d_writedata[16]~reg0_q ),
	.d_writedata_27(\nios2_qsys_0|d_writedata[27]~reg0_q ),
	.d_writedata_19(\nios2_qsys_0|d_writedata[19]~reg0_q ),
	.d_writedata_26(\nios2_qsys_0|d_writedata[26]~reg0_q ),
	.d_writedata_18(\nios2_qsys_0|d_writedata[18]~reg0_q ),
	.d_writedata_23(\nios2_qsys_0|d_writedata[23]~reg0_q ),
	.d_writedata_15(\nios2_qsys_0|d_writedata[15]~reg0_q ),
	.d_writedata_22(\nios2_qsys_0|d_writedata[22]~reg0_q ),
	.d_writedata_14(\nios2_qsys_0|d_writedata[14]~reg0_q ),
	.d_byteenable_1(\nios2_qsys_0|d_byteenable[1]~reg0_q ),
	.d_writedata_2(\nios2_qsys_0|d_writedata[2]~reg0_q ),
	.d_writedata_0(\nios2_qsys_0|d_writedata[0]~reg0_q ),
	.d_writedata_3(\nios2_qsys_0|d_writedata[3]~reg0_q ),
	.d_writedata_1(\nios2_qsys_0|d_writedata[1]~reg0_q ),
	.d_writedata_6(\nios2_qsys_0|d_writedata[6]~reg0_q ),
	.d_writedata_4(\nios2_qsys_0|d_writedata[4]~reg0_q ),
	.d_writedata_7(\nios2_qsys_0|d_writedata[7]~reg0_q ),
	.d_writedata_5(\nios2_qsys_0|d_writedata[5]~reg0_q ),
	.clk_clk(\clk_clk~input_o ));

embedded_system_embedded_system_nios2_qsys_0 nios2_qsys_0(
	.readdata_2(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[2]~q ),
	.readdata_10(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[10]~q ),
	.readdata_18(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[18]~q ),
	.readdata_26(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[26]~q ),
	.readdata_7(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[7]~q ),
	.readdata_23(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[23]~q ),
	.readdata_15(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[15]~q ),
	.readdata_31(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[31]~q ),
	.readdata_29(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[29]~q ),
	.readdata_13(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[13]~q ),
	.readdata_28(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[28]~q ),
	.readdata_12(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[12]~q ),
	.readdata_27(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[27]~q ),
	.readdata_11(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[11]~q ),
	.readdata_25(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[25]~q ),
	.readdata_9(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[9]~q ),
	.readdata_24(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[24]~q ),
	.readdata_8(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[8]~q ),
	.readdata_6(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[6]~q ),
	.readdata_14(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[14]~q ),
	.readdata_22(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[22]~q ),
	.readdata_30(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[30]~q ),
	.readdata_5(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[5]~q ),
	.readdata_21(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[21]~q ),
	.readdata_4(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[4]~q ),
	.readdata_20(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[20]~q ),
	.readdata_3(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[3]~q ),
	.readdata_19(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[19]~q ),
	.readdata_1(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[1]~q ),
	.readdata_17(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[17]~q ),
	.readdata_0(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[0]~q ),
	.readdata_16(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[16]~q ),
	.sr_0(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[0]~q ),
	.ir_out_0(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[0]~q ),
	.ir_out_1(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[1]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.hold_waitrequest(\mm_interconnect_0|nios2_qsys_0_data_master_agent|hold_waitrequest~q ),
	.d_address_offset_field_0(\nios2_qsys_0|d_address_offset_field[0]~q ),
	.d_write(\nios2_qsys_0|d_write~reg0_q ),
	.d_address_tag_field_2(\nios2_qsys_0|d_address_tag_field[2]~q ),
	.d_address_tag_field_1(\nios2_qsys_0|d_address_tag_field[1]~q ),
	.d_address_tag_field_0(\nios2_qsys_0|d_address_tag_field[0]~q ),
	.d_address_line_field_5(\nios2_qsys_0|d_address_line_field[5]~q ),
	.d_address_line_field_4(\nios2_qsys_0|d_address_line_field[4]~q ),
	.d_address_line_field_3(\nios2_qsys_0|d_address_line_field[3]~q ),
	.d_address_line_field_2(\nios2_qsys_0|d_address_line_field[2]~q ),
	.d_address_line_field_1(\nios2_qsys_0|d_address_line_field[1]~q ),
	.d_address_line_field_0(\nios2_qsys_0|d_address_line_field[0]~q ),
	.d_address_offset_field_2(\nios2_qsys_0|d_address_offset_field[2]~q ),
	.d_address_offset_field_1(\nios2_qsys_0|d_address_offset_field[1]~q ),
	.d_writedata_11(\nios2_qsys_0|d_writedata[11]~reg0_q ),
	.d_byteenable_0(\nios2_qsys_0|d_byteenable[0]~reg0_q ),
	.d_writedata_10(\nios2_qsys_0|d_writedata[10]~reg0_q ),
	.d_writedata_9(\nios2_qsys_0|d_writedata[9]~reg0_q ),
	.d_writedata_8(\nios2_qsys_0|d_writedata[8]~reg0_q ),
	.d_writedata_13(\nios2_qsys_0|d_writedata[13]~reg0_q ),
	.d_writedata_12(\nios2_qsys_0|d_writedata[12]~reg0_q ),
	.d_writedata_21(\nios2_qsys_0|d_writedata[21]~reg0_q ),
	.d_writedata_20(\nios2_qsys_0|d_writedata[20]~reg0_q ),
	.d_writedata_25(\nios2_qsys_0|d_writedata[25]~reg0_q ),
	.d_writedata_17(\nios2_qsys_0|d_writedata[17]~reg0_q ),
	.d_writedata_24(\nios2_qsys_0|d_writedata[24]~reg0_q ),
	.d_writedata_16(\nios2_qsys_0|d_writedata[16]~reg0_q ),
	.d_writedata_27(\nios2_qsys_0|d_writedata[27]~reg0_q ),
	.d_writedata_19(\nios2_qsys_0|d_writedata[19]~reg0_q ),
	.d_writedata_26(\nios2_qsys_0|d_writedata[26]~reg0_q ),
	.d_writedata_18(\nios2_qsys_0|d_writedata[18]~reg0_q ),
	.d_writedata_23(\nios2_qsys_0|d_writedata[23]~reg0_q ),
	.d_writedata_15(\nios2_qsys_0|d_writedata[15]~reg0_q ),
	.d_writedata_22(\nios2_qsys_0|d_writedata[22]~reg0_q ),
	.d_writedata_14(\nios2_qsys_0|d_writedata[14]~reg0_q ),
	.d_read(\nios2_qsys_0|d_read~reg0_q ),
	.suppress_change_dest_id(\mm_interconnect_0|nios2_qsys_0_data_master_limiter|suppress_change_dest_id~0_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ),
	.jtag_debug_module_waitrequest(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\mm_interconnect_0|cmd_demux|WideOr0~combout ),
	.av_waitrequest(\mm_interconnect_0|nios2_qsys_0_data_master_agent|av_waitrequest~combout ),
	.d_byteenable_1(\nios2_qsys_0|d_byteenable[1]~reg0_q ),
	.d_writedata_2(\nios2_qsys_0|d_writedata[2]~reg0_q ),
	.d_writedata_0(\nios2_qsys_0|d_writedata[0]~reg0_q ),
	.d_writedata_3(\nios2_qsys_0|d_writedata[3]~reg0_q ),
	.d_writedata_1(\nios2_qsys_0|d_writedata[1]~reg0_q ),
	.hbreak_enabled1(\nios2_qsys_0|hbreak_enabled~q ),
	.i_read(\nios2_qsys_0|i_read~reg0_q ),
	.src0_valid(\mm_interconnect_0|cmd_demux_001|src0_valid~0_combout ),
	.ic_fill_tag_1(\nios2_qsys_0|ic_fill_tag[1]~q ),
	.ic_fill_tag_0(\nios2_qsys_0|ic_fill_tag[0]~q ),
	.ic_fill_line_6(\nios2_qsys_0|ic_fill_line[6]~q ),
	.Equal1(\mm_interconnect_0|router_001|Equal1~0_combout ),
	.src0_valid1(\mm_interconnect_0|cmd_demux_001|src0_valid~1_combout ),
	.src1_valid(\mm_interconnect_0|cmd_demux|src1_valid~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_001|saved_grant[1]~q ),
	.rf_source_valid(\mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent|rf_source_valid~0_combout ),
	.d_writedata_6(\nios2_qsys_0|d_writedata[6]~reg0_q ),
	.d_writedata_4(\nios2_qsys_0|d_writedata[4]~reg0_q ),
	.d_writedata_7(\nios2_qsys_0|d_writedata[7]~reg0_q ),
	.d_writedata_5(\nios2_qsys_0|d_writedata[5]~reg0_q ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.d_readdatavalid(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.suppress_change_dest_id1(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|suppress_change_dest_id~0_combout ),
	.WideOr01(\mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ),
	.WideOr02(\mm_interconnect_0|cmd_demux_001|WideOr0~1_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|nonposted_cmd_accepted~combout ),
	.ic_fill_line_5(\nios2_qsys_0|ic_fill_line[5]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_001|src_data[46]~combout ),
	.src_payload(\mm_interconnect_0|cmd_mux_001|src_payload~0_combout ),
	.ic_fill_ap_offset_0(\nios2_qsys_0|ic_fill_ap_offset[0]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_001|src_data[38]~combout ),
	.ic_fill_line_1(\nios2_qsys_0|ic_fill_line[1]~q ),
	.src_data_42(\mm_interconnect_0|cmd_mux_001|src_data[42]~combout ),
	.ic_fill_line_0(\nios2_qsys_0|ic_fill_line[0]~q ),
	.src_data_41(\mm_interconnect_0|cmd_mux_001|src_data[41]~combout ),
	.ic_fill_ap_offset_2(\nios2_qsys_0|ic_fill_ap_offset[2]~q ),
	.src_data_40(\mm_interconnect_0|cmd_mux_001|src_data[40]~combout ),
	.ic_fill_ap_offset_1(\nios2_qsys_0|ic_fill_ap_offset[1]~q ),
	.src_data_39(\mm_interconnect_0|cmd_mux_001|src_data[39]~combout ),
	.ic_fill_line_4(\nios2_qsys_0|ic_fill_line[4]~q ),
	.src_data_45(\mm_interconnect_0|cmd_mux_001|src_data[45]~combout ),
	.ic_fill_line_3(\nios2_qsys_0|ic_fill_line[3]~q ),
	.src_data_44(\mm_interconnect_0|cmd_mux_001|src_data[44]~combout ),
	.ic_fill_line_2(\nios2_qsys_0|ic_fill_line[2]~q ),
	.src_data_43(\mm_interconnect_0|cmd_mux_001|src_data[43]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_001|src_payload~1_combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_001|src_data[32]~combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_001|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_001|src_payload~3_combout ),
	.WideOr1(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.d_readdata({\mm_interconnect_0|rsp_mux|src_data[31]~combout ,\mm_interconnect_0|rsp_mux|src_data[30]~combout ,\mm_interconnect_0|rsp_mux|src_data[29]~combout ,\mm_interconnect_0|rsp_mux|src_data[28]~combout ,\mm_interconnect_0|rsp_mux|src_data[27]~combout ,
\mm_interconnect_0|rsp_mux|src_data[26]~combout ,\mm_interconnect_0|rsp_mux|src_data[25]~combout ,\mm_interconnect_0|rsp_mux|src_data[24]~combout ,\mm_interconnect_0|rsp_mux|src_data[23]~combout ,\mm_interconnect_0|rsp_mux|src_data[22]~combout ,
\mm_interconnect_0|rsp_mux|src_data[21]~combout ,\mm_interconnect_0|rsp_mux|src_data[20]~combout ,\mm_interconnect_0|rsp_mux|src_data[19]~combout ,\mm_interconnect_0|rsp_mux|src_data[18]~combout ,\mm_interconnect_0|rsp_mux|src_data[17]~combout ,
\mm_interconnect_0|rsp_mux|src_data[16]~combout ,\mm_interconnect_0|rsp_mux|src_data[15]~combout ,\mm_interconnect_0|rsp_mux|src_data[14]~combout ,\mm_interconnect_0|rsp_mux|src_data[13]~combout ,\mm_interconnect_0|rsp_mux|src_data[12]~combout ,
\mm_interconnect_0|rsp_mux|src_data[11]~combout ,\mm_interconnect_0|rsp_mux|src_data[10]~combout ,\mm_interconnect_0|rsp_mux|src_data[9]~combout ,\mm_interconnect_0|rsp_mux|src_data[8]~combout ,\mm_interconnect_0|rsp_mux|src_data[7]~combout ,
\mm_interconnect_0|rsp_mux|src_data[6]~combout ,\mm_interconnect_0|rsp_mux|src_data[5]~combout ,\mm_interconnect_0|rsp_mux|src_data[4]~combout ,\mm_interconnect_0|rsp_mux|src_data[3]~combout ,\mm_interconnect_0|rsp_mux|src_data[2]~combout ,
\mm_interconnect_0|rsp_mux|src_data[1]~combout ,\mm_interconnect_0|rsp_mux|src_data[0]~combout }),
	.jtag_debug_module_resetrequest(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_oci_debug|resetrequest~q ),
	.src_payload4(\mm_interconnect_0|cmd_mux_001|src_payload~4_combout ),
	.i_readdata({\mm_interconnect_0|rsp_mux_001|src_data[31]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[30]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[29]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[28]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[27]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[26]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[25]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[24]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[23]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[22]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[21]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[20]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[19]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[18]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[17]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[16]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[15]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[14]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[13]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[12]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[11]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[10]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[9]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[8]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[7]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[6]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[5]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[4]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[3]~combout ,
\mm_interconnect_0|rsp_mux_001|src_data[2]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[1]~combout ,\mm_interconnect_0|rsp_mux_001|src_data[0]~combout }),
	.d_byteenable_2(\nios2_qsys_0|d_byteenable[2]~reg0_q ),
	.d_byteenable_3(\nios2_qsys_0|d_byteenable[3]~reg0_q ),
	.d_writedata_31(\nios2_qsys_0|d_writedata[31]~reg0_q ),
	.d_writedata_29(\nios2_qsys_0|d_writedata[29]~reg0_q ),
	.d_writedata_28(\nios2_qsys_0|d_writedata[28]~reg0_q ),
	.d_writedata_30(\nios2_qsys_0|d_writedata[30]~reg0_q ),
	.src_payload5(\mm_interconnect_0|cmd_mux_001|src_payload~5_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_001|src_data[35]~combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_001|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_001|src_payload~7_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_001|src_data[34]~combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_001|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_001|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_001|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_001|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_001|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_001|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_001|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_001|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_001|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_001|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_001|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_001|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_001|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_001|src_payload~21_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_001|src_data[33]~combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_001|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_001|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_001|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_001|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_001|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_001|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_001|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_001|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_001|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_001|src_payload~31_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_001|src_payload~32_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TCKUTAP ),
	.altera_internal_jtag1(\altera_internal_jtag~TDIUTAP ),
	.NJQG9082(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.state_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.state_4(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.splitter_nodes_receive_0_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.virtual_ir_scan_reg(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.state_8(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.irf_reg_0_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.clk_clk(\clk_clk~input_o ));

embedded_system_embedded_system_mm_interconnect_0 mm_interconnect_0(
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.readdata_2(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[2]~q ),
	.readdata_10(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[10]~q ),
	.readdata_18(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[18]~q ),
	.readdata_26(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[26]~q ),
	.readdata_7(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[7]~q ),
	.readdata_23(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[23]~q ),
	.readdata_15(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[15]~q ),
	.readdata_31(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[31]~q ),
	.readdata_29(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[29]~q ),
	.readdata_13(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[13]~q ),
	.readdata_28(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[28]~q ),
	.readdata_12(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[12]~q ),
	.readdata_27(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[27]~q ),
	.readdata_11(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[11]~q ),
	.readdata_25(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[25]~q ),
	.readdata_9(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[9]~q ),
	.readdata_24(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[24]~q ),
	.readdata_8(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[8]~q ),
	.readdata_6(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[6]~q ),
	.readdata_14(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[14]~q ),
	.readdata_22(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[22]~q ),
	.readdata_30(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[30]~q ),
	.readdata_5(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[5]~q ),
	.readdata_21(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[21]~q ),
	.readdata_4(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[4]~q ),
	.readdata_20(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[20]~q ),
	.readdata_3(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[3]~q ),
	.readdata_19(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[19]~q ),
	.readdata_1(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[1]~q ),
	.readdata_17(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[17]~q ),
	.readdata_0(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[0]~q ),
	.readdata_16(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|readdata[16]~q ),
	.r_sync_rst(\rst_controller|r_sync_rst~q ),
	.wait_latency_counter_1(\mm_interconnect_0|ad9833_comp_0_avalon_slave_0_translator|wait_latency_counter[1]~q ),
	.wait_latency_counter_0(\mm_interconnect_0|ad9833_comp_0_avalon_slave_0_translator|wait_latency_counter[0]~q ),
	.hold_waitrequest(\mm_interconnect_0|nios2_qsys_0_data_master_agent|hold_waitrequest~q ),
	.d_address_offset_field_0(\nios2_qsys_0|d_address_offset_field[0]~q ),
	.d_write(\nios2_qsys_0|d_write~reg0_q ),
	.d_address_tag_field_2(\nios2_qsys_0|d_address_tag_field[2]~q ),
	.d_address_tag_field_1(\nios2_qsys_0|d_address_tag_field[1]~q ),
	.d_address_tag_field_0(\nios2_qsys_0|d_address_tag_field[0]~q ),
	.d_address_line_field_5(\nios2_qsys_0|d_address_line_field[5]~q ),
	.d_address_line_field_4(\nios2_qsys_0|d_address_line_field[4]~q ),
	.d_address_line_field_3(\nios2_qsys_0|d_address_line_field[3]~q ),
	.d_address_line_field_2(\nios2_qsys_0|d_address_line_field[2]~q ),
	.d_address_line_field_1(\nios2_qsys_0|d_address_line_field[1]~q ),
	.d_address_line_field_0(\nios2_qsys_0|d_address_line_field[0]~q ),
	.d_address_offset_field_2(\nios2_qsys_0|d_address_offset_field[2]~q ),
	.d_address_offset_field_1(\nios2_qsys_0|d_address_offset_field[1]~q ),
	.m0_write(\mm_interconnect_0|ad9833_comp_0_avalon_slave_0_agent|m0_write~0_combout ),
	.d_writedata_11(\nios2_qsys_0|d_writedata[11]~reg0_q ),
	.d_byteenable_0(\nios2_qsys_0|d_byteenable[0]~reg0_q ),
	.d_writedata_10(\nios2_qsys_0|d_writedata[10]~reg0_q ),
	.d_writedata_9(\nios2_qsys_0|d_writedata[9]~reg0_q ),
	.d_writedata_8(\nios2_qsys_0|d_writedata[8]~reg0_q ),
	.d_writedata_13(\nios2_qsys_0|d_writedata[13]~reg0_q ),
	.d_writedata_12(\nios2_qsys_0|d_writedata[12]~reg0_q ),
	.d_writedata_21(\nios2_qsys_0|d_writedata[21]~reg0_q ),
	.d_writedata_20(\nios2_qsys_0|d_writedata[20]~reg0_q ),
	.d_writedata_25(\nios2_qsys_0|d_writedata[25]~reg0_q ),
	.d_writedata_17(\nios2_qsys_0|d_writedata[17]~reg0_q ),
	.d_writedata_24(\nios2_qsys_0|d_writedata[24]~reg0_q ),
	.d_writedata_16(\nios2_qsys_0|d_writedata[16]~reg0_q ),
	.d_writedata_27(\nios2_qsys_0|d_writedata[27]~reg0_q ),
	.d_writedata_19(\nios2_qsys_0|d_writedata[19]~reg0_q ),
	.d_writedata_26(\nios2_qsys_0|d_writedata[26]~reg0_q ),
	.d_writedata_18(\nios2_qsys_0|d_writedata[18]~reg0_q ),
	.d_writedata_23(\nios2_qsys_0|d_writedata[23]~reg0_q ),
	.d_writedata_15(\nios2_qsys_0|d_writedata[15]~reg0_q ),
	.d_writedata_22(\nios2_qsys_0|d_writedata[22]~reg0_q ),
	.d_writedata_14(\nios2_qsys_0|d_writedata[14]~reg0_q ),
	.d_read(\nios2_qsys_0|d_read~reg0_q ),
	.suppress_change_dest_id(\mm_interconnect_0|nios2_qsys_0_data_master_limiter|suppress_change_dest_id~0_combout ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_001|saved_grant[0]~q ),
	.waitrequest(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_ocimem|waitrequest~q ),
	.mem_used_1(\mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem_used[1]~q ),
	.saved_grant_01(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.mem_used_11(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.WideOr0(\mm_interconnect_0|cmd_demux|WideOr0~combout ),
	.av_waitrequest(\mm_interconnect_0|nios2_qsys_0_data_master_agent|av_waitrequest~combout ),
	.d_byteenable_1(\nios2_qsys_0|d_byteenable[1]~reg0_q ),
	.d_writedata_2(\nios2_qsys_0|d_writedata[2]~reg0_q ),
	.d_writedata_0(\nios2_qsys_0|d_writedata[0]~reg0_q ),
	.d_writedata_3(\nios2_qsys_0|d_writedata[3]~reg0_q ),
	.d_writedata_1(\nios2_qsys_0|d_writedata[1]~reg0_q ),
	.hbreak_enabled(\nios2_qsys_0|hbreak_enabled~q ),
	.i_read(\nios2_qsys_0|i_read~reg0_q ),
	.src0_valid(\mm_interconnect_0|cmd_demux_001|src0_valid~0_combout ),
	.ic_fill_tag_1(\nios2_qsys_0|ic_fill_tag[1]~q ),
	.ic_fill_tag_0(\nios2_qsys_0|ic_fill_tag[0]~q ),
	.ic_fill_line_6(\nios2_qsys_0|ic_fill_line[6]~q ),
	.Equal1(\mm_interconnect_0|router_001|Equal1~0_combout ),
	.src0_valid1(\mm_interconnect_0|cmd_demux_001|src0_valid~1_combout ),
	.src1_valid(\mm_interconnect_0|cmd_demux|src1_valid~0_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_001|saved_grant[1]~q ),
	.rf_source_valid(\mm_interconnect_0|nios2_qsys_0_jtag_debug_module_agent|rf_source_valid~0_combout ),
	.src1_valid1(\mm_interconnect_0|cmd_demux_001|src1_valid~0_combout ),
	.src2_valid(\mm_interconnect_0|cmd_demux|src2_valid~2_combout ),
	.saved_grant_11(\mm_interconnect_0|cmd_mux_002|saved_grant[1]~q ),
	.d_writedata_6(\nios2_qsys_0|d_writedata[6]~reg0_q ),
	.d_writedata_4(\nios2_qsys_0|d_writedata[4]~reg0_q ),
	.d_writedata_7(\nios2_qsys_0|d_writedata[7]~reg0_q ),
	.d_writedata_5(\nios2_qsys_0|d_writedata[5]~reg0_q ),
	.WideOr1(\mm_interconnect_0|rsp_mux|WideOr1~combout ),
	.suppress_change_dest_id1(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|suppress_change_dest_id~0_combout ),
	.WideOr01(\mm_interconnect_0|cmd_demux_001|WideOr0~0_combout ),
	.WideOr02(\mm_interconnect_0|cmd_demux_001|WideOr0~1_combout ),
	.nonposted_cmd_accepted(\mm_interconnect_0|nios2_qsys_0_instruction_master_limiter|nonposted_cmd_accepted~combout ),
	.ic_fill_line_5(\nios2_qsys_0|ic_fill_line[5]~q ),
	.src_data_46(\mm_interconnect_0|cmd_mux_001|src_data[46]~combout ),
	.src_payload(\mm_interconnect_0|cmd_mux_001|src_payload~0_combout ),
	.ic_fill_ap_offset_0(\nios2_qsys_0|ic_fill_ap_offset[0]~q ),
	.src_data_38(\mm_interconnect_0|cmd_mux_001|src_data[38]~combout ),
	.ic_fill_line_1(\nios2_qsys_0|ic_fill_line[1]~q ),
	.src_data_42(\mm_interconnect_0|cmd_mux_001|src_data[42]~combout ),
	.ic_fill_line_0(\nios2_qsys_0|ic_fill_line[0]~q ),
	.src_data_41(\mm_interconnect_0|cmd_mux_001|src_data[41]~combout ),
	.ic_fill_ap_offset_2(\nios2_qsys_0|ic_fill_ap_offset[2]~q ),
	.src_data_40(\mm_interconnect_0|cmd_mux_001|src_data[40]~combout ),
	.ic_fill_ap_offset_1(\nios2_qsys_0|ic_fill_ap_offset[1]~q ),
	.src_data_39(\mm_interconnect_0|cmd_mux_001|src_data[39]~combout ),
	.ic_fill_line_4(\nios2_qsys_0|ic_fill_line[4]~q ),
	.src_data_45(\mm_interconnect_0|cmd_mux_001|src_data[45]~combout ),
	.ic_fill_line_3(\nios2_qsys_0|ic_fill_line[3]~q ),
	.src_data_44(\mm_interconnect_0|cmd_mux_001|src_data[44]~combout ),
	.ic_fill_line_2(\nios2_qsys_0|ic_fill_line[2]~q ),
	.src_data_43(\mm_interconnect_0|cmd_mux_001|src_data[43]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_001|src_payload~1_combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_001|src_data[32]~combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_001|src_payload~2_combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_001|src_payload~3_combout ),
	.WideOr11(\mm_interconnect_0|rsp_mux_001|WideOr1~combout ),
	.src_data_2(\mm_interconnect_0|rsp_mux|src_data[2]~combout ),
	.src_data_10(\mm_interconnect_0|rsp_mux|src_data[10]~combout ),
	.src_data_18(\mm_interconnect_0|rsp_mux|src_data[18]~combout ),
	.src_data_26(\mm_interconnect_0|rsp_mux|src_data[26]~combout ),
	.src_data_7(\mm_interconnect_0|rsp_mux|src_data[7]~combout ),
	.src_data_23(\mm_interconnect_0|rsp_mux|src_data[23]~combout ),
	.src_data_15(\mm_interconnect_0|rsp_mux|src_data[15]~combout ),
	.src_data_31(\mm_interconnect_0|rsp_mux|src_data[31]~combout ),
	.src_data_29(\mm_interconnect_0|rsp_mux|src_data[29]~combout ),
	.src_data_13(\mm_interconnect_0|rsp_mux|src_data[13]~combout ),
	.src_data_28(\mm_interconnect_0|rsp_mux|src_data[28]~combout ),
	.src_data_12(\mm_interconnect_0|rsp_mux|src_data[12]~combout ),
	.src_data_27(\mm_interconnect_0|rsp_mux|src_data[27]~combout ),
	.src_data_11(\mm_interconnect_0|rsp_mux|src_data[11]~combout ),
	.src_data_25(\mm_interconnect_0|rsp_mux|src_data[25]~combout ),
	.src_data_9(\mm_interconnect_0|rsp_mux|src_data[9]~combout ),
	.src_data_24(\mm_interconnect_0|rsp_mux|src_data[24]~combout ),
	.src_data_8(\mm_interconnect_0|rsp_mux|src_data[8]~combout ),
	.src_data_6(\mm_interconnect_0|rsp_mux|src_data[6]~combout ),
	.src_data_14(\mm_interconnect_0|rsp_mux|src_data[14]~combout ),
	.src_data_22(\mm_interconnect_0|rsp_mux|src_data[22]~combout ),
	.src_data_30(\mm_interconnect_0|rsp_mux|src_data[30]~combout ),
	.src_data_5(\mm_interconnect_0|rsp_mux|src_data[5]~combout ),
	.src_data_21(\mm_interconnect_0|rsp_mux|src_data[21]~combout ),
	.src_data_4(\mm_interconnect_0|rsp_mux|src_data[4]~combout ),
	.src_data_20(\mm_interconnect_0|rsp_mux|src_data[20]~combout ),
	.src_data_3(\mm_interconnect_0|rsp_mux|src_data[3]~combout ),
	.src_data_19(\mm_interconnect_0|rsp_mux|src_data[19]~combout ),
	.src_data_1(\mm_interconnect_0|rsp_mux|src_data[1]~combout ),
	.src_data_17(\mm_interconnect_0|rsp_mux|src_data[17]~combout ),
	.src_data_0(\mm_interconnect_0|rsp_mux|src_data[0]~combout ),
	.src_data_16(\mm_interconnect_0|rsp_mux|src_data[16]~combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_001|src_payload~4_combout ),
	.src_data_51(\mm_interconnect_0|rsp_mux_001|src_data[5]~combout ),
	.src_data_33(\mm_interconnect_0|rsp_mux_001|src_data[3]~combout ),
	.src_data_110(\mm_interconnect_0|rsp_mux_001|src_data[1]~combout ),
	.src_data_47(\mm_interconnect_0|rsp_mux_001|src_data[4]~combout ),
	.src_data_210(\mm_interconnect_0|rsp_mux_001|src_data[2]~combout ),
	.src_data_281(\mm_interconnect_0|rsp_mux_001|src_data[28]~combout ),
	.src_data_311(\mm_interconnect_0|rsp_mux_001|src_data[31]~combout ),
	.src_data_271(\mm_interconnect_0|rsp_mux_001|src_data[27]~combout ),
	.src_data_291(\mm_interconnect_0|rsp_mux_001|src_data[29]~combout ),
	.src_data_301(\mm_interconnect_0|rsp_mux_001|src_data[30]~combout ),
	.src_data_01(\mm_interconnect_0|rsp_mux_001|src_data[0]~combout ),
	.src_data_231(\mm_interconnect_0|rsp_mux_001|src_data[23]~combout ),
	.src_data_261(\mm_interconnect_0|rsp_mux_001|src_data[26]~combout ),
	.src_data_221(\mm_interconnect_0|rsp_mux_001|src_data[22]~combout ),
	.src_data_241(\mm_interconnect_0|rsp_mux_001|src_data[24]~combout ),
	.src_data_251(\mm_interconnect_0|rsp_mux_001|src_data[25]~combout ),
	.src_data_161(\mm_interconnect_0|rsp_mux_001|src_data[16]~combout ),
	.src_data_151(\mm_interconnect_0|rsp_mux_001|src_data[15]~combout ),
	.src_data_131(\mm_interconnect_0|rsp_mux_001|src_data[13]~combout ),
	.src_data_141(\mm_interconnect_0|rsp_mux_001|src_data[14]~combout ),
	.src_data_121(\mm_interconnect_0|rsp_mux_001|src_data[12]~combout ),
	.src_data_111(\mm_interconnect_0|rsp_mux_001|src_data[11]~combout ),
	.src_data_81(\mm_interconnect_0|rsp_mux_001|src_data[8]~combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_data_381(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_391(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_401(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_411(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_421(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_data_431(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_441(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_451(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_461(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.src_data_471(\mm_interconnect_0|cmd_mux_002|src_data[47]~combout ),
	.src_data_321(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.src_data_331(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.d_byteenable_2(\nios2_qsys_0|d_byteenable[2]~reg0_q ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.d_byteenable_3(\nios2_qsys_0|d_byteenable[3]~reg0_q ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_data_191(\mm_interconnect_0|rsp_mux_001|src_data[19]~combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.d_writedata_31(\nios2_qsys_0|d_writedata[31]~reg0_q ),
	.src_payload12(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.d_writedata_29(\nios2_qsys_0|d_writedata[29]~reg0_q ),
	.src_payload13(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_data_181(\mm_interconnect_0|rsp_mux_001|src_data[18]~combout ),
	.d_writedata_28(\nios2_qsys_0|d_writedata[28]~reg0_q ),
	.src_payload15(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_data_171(\mm_interconnect_0|rsp_mux_001|src_data[17]~combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.d_writedata_30(\nios2_qsys_0|d_writedata[30]~reg0_q ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_data_101(\mm_interconnect_0|rsp_mux_001|src_data[10]~combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_data_91(\mm_interconnect_0|rsp_mux_001|src_data[9]~combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload32(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload33(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload34(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload35(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload36(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.src_data_211(\mm_interconnect_0|rsp_mux_001|src_data[21]~combout ),
	.src_data_201(\mm_interconnect_0|rsp_mux_001|src_data[20]~combout ),
	.src_data_71(\mm_interconnect_0|rsp_mux_001|src_data[7]~combout ),
	.src_data_61(\mm_interconnect_0|rsp_mux_001|src_data[6]~combout ),
	.src_payload37(\mm_interconnect_0|cmd_mux_001|src_payload~5_combout ),
	.src_data_351(\mm_interconnect_0|cmd_mux_001|src_data[35]~combout ),
	.src_payload38(\mm_interconnect_0|cmd_mux_001|src_payload~6_combout ),
	.src_payload39(\mm_interconnect_0|cmd_mux_001|src_payload~7_combout ),
	.src_data_341(\mm_interconnect_0|cmd_mux_001|src_data[34]~combout ),
	.src_payload40(\mm_interconnect_0|cmd_mux_001|src_payload~8_combout ),
	.src_payload41(\mm_interconnect_0|cmd_mux_001|src_payload~9_combout ),
	.src_payload42(\mm_interconnect_0|cmd_mux_001|src_payload~10_combout ),
	.src_payload43(\mm_interconnect_0|cmd_mux_001|src_payload~11_combout ),
	.src_payload44(\mm_interconnect_0|cmd_mux_001|src_payload~12_combout ),
	.src_payload45(\mm_interconnect_0|cmd_mux_001|src_payload~13_combout ),
	.src_payload46(\mm_interconnect_0|cmd_mux_001|src_payload~14_combout ),
	.src_payload47(\mm_interconnect_0|cmd_mux_001|src_payload~15_combout ),
	.src_payload48(\mm_interconnect_0|cmd_mux_001|src_payload~16_combout ),
	.src_payload49(\mm_interconnect_0|cmd_mux_001|src_payload~17_combout ),
	.src_payload50(\mm_interconnect_0|cmd_mux_001|src_payload~18_combout ),
	.src_payload51(\mm_interconnect_0|cmd_mux_001|src_payload~19_combout ),
	.src_payload52(\mm_interconnect_0|cmd_mux_001|src_payload~20_combout ),
	.src_payload53(\mm_interconnect_0|cmd_mux_001|src_payload~21_combout ),
	.src_data_332(\mm_interconnect_0|cmd_mux_001|src_data[33]~combout ),
	.src_payload54(\mm_interconnect_0|cmd_mux_001|src_payload~22_combout ),
	.src_payload55(\mm_interconnect_0|cmd_mux_001|src_payload~23_combout ),
	.src_payload56(\mm_interconnect_0|cmd_mux_001|src_payload~24_combout ),
	.src_payload57(\mm_interconnect_0|cmd_mux_001|src_payload~25_combout ),
	.src_payload58(\mm_interconnect_0|cmd_mux_001|src_payload~26_combout ),
	.src_payload59(\mm_interconnect_0|cmd_mux_001|src_payload~27_combout ),
	.src_payload60(\mm_interconnect_0|cmd_mux_001|src_payload~28_combout ),
	.src_payload61(\mm_interconnect_0|cmd_mux_001|src_payload~29_combout ),
	.src_payload62(\mm_interconnect_0|cmd_mux_001|src_payload~30_combout ),
	.src_payload63(\mm_interconnect_0|cmd_mux_001|src_payload~31_combout ),
	.src_payload64(\mm_interconnect_0|cmd_mux_001|src_payload~32_combout ),
	.clk_clk(\clk_clk~input_o ));

embedded_system_embedded_system_onchip_memory2_0 onchip_memory2_0(
	.q_a_2(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[2] ),
	.q_a_10(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_18(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_26(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_7(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_23(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_15(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_31(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[31] ),
	.q_a_29(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_13(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_28(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_12(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_27(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_11(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_25(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[25] ),
	.q_a_9(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_24(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_8(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_6(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_14(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_22(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[22] ),
	.q_a_30(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_5(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_21(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_4(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[4] ),
	.q_a_20(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_3(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[3] ),
	.q_a_19(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[19] ),
	.q_a_1(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_17(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_0(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_16(\onchip_memory2_0|the_altsyncram|auto_generated|q_a[16] ),
	.d_write(\nios2_qsys_0|d_write~reg0_q ),
	.saved_grant_0(\mm_interconnect_0|cmd_mux_002|saved_grant[0]~q ),
	.mem_used_1(\mm_interconnect_0|onchip_memory2_0_s1_agent_rsp_fifo|mem_used[1]~q ),
	.src1_valid(\mm_interconnect_0|cmd_demux_001|src1_valid~0_combout ),
	.src2_valid(\mm_interconnect_0|cmd_demux|src2_valid~2_combout ),
	.saved_grant_1(\mm_interconnect_0|cmd_mux_002|saved_grant[1]~q ),
	.r_early_rst(\rst_controller|r_early_rst~q ),
	.src_payload(\mm_interconnect_0|cmd_mux_002|src_payload~0_combout ),
	.src_data_38(\mm_interconnect_0|cmd_mux_002|src_data[38]~combout ),
	.src_data_39(\mm_interconnect_0|cmd_mux_002|src_data[39]~combout ),
	.src_data_40(\mm_interconnect_0|cmd_mux_002|src_data[40]~combout ),
	.src_data_41(\mm_interconnect_0|cmd_mux_002|src_data[41]~combout ),
	.src_data_42(\mm_interconnect_0|cmd_mux_002|src_data[42]~combout ),
	.src_data_43(\mm_interconnect_0|cmd_mux_002|src_data[43]~combout ),
	.src_data_44(\mm_interconnect_0|cmd_mux_002|src_data[44]~combout ),
	.src_data_45(\mm_interconnect_0|cmd_mux_002|src_data[45]~combout ),
	.src_data_46(\mm_interconnect_0|cmd_mux_002|src_data[46]~combout ),
	.src_data_47(\mm_interconnect_0|cmd_mux_002|src_data[47]~combout ),
	.src_data_32(\mm_interconnect_0|cmd_mux_002|src_data[32]~combout ),
	.src_payload1(\mm_interconnect_0|cmd_mux_002|src_payload~1_combout ),
	.src_data_33(\mm_interconnect_0|cmd_mux_002|src_data[33]~combout ),
	.src_payload2(\mm_interconnect_0|cmd_mux_002|src_payload~2_combout ),
	.src_data_34(\mm_interconnect_0|cmd_mux_002|src_data[34]~combout ),
	.src_payload3(\mm_interconnect_0|cmd_mux_002|src_payload~3_combout ),
	.src_data_35(\mm_interconnect_0|cmd_mux_002|src_data[35]~combout ),
	.src_payload4(\mm_interconnect_0|cmd_mux_002|src_payload~4_combout ),
	.src_payload5(\mm_interconnect_0|cmd_mux_002|src_payload~5_combout ),
	.src_payload6(\mm_interconnect_0|cmd_mux_002|src_payload~6_combout ),
	.src_payload7(\mm_interconnect_0|cmd_mux_002|src_payload~7_combout ),
	.src_payload8(\mm_interconnect_0|cmd_mux_002|src_payload~8_combout ),
	.src_payload9(\mm_interconnect_0|cmd_mux_002|src_payload~9_combout ),
	.src_payload10(\mm_interconnect_0|cmd_mux_002|src_payload~10_combout ),
	.src_payload11(\mm_interconnect_0|cmd_mux_002|src_payload~11_combout ),
	.src_payload12(\mm_interconnect_0|cmd_mux_002|src_payload~12_combout ),
	.src_payload13(\mm_interconnect_0|cmd_mux_002|src_payload~13_combout ),
	.src_payload14(\mm_interconnect_0|cmd_mux_002|src_payload~14_combout ),
	.src_payload15(\mm_interconnect_0|cmd_mux_002|src_payload~15_combout ),
	.src_payload16(\mm_interconnect_0|cmd_mux_002|src_payload~16_combout ),
	.src_payload17(\mm_interconnect_0|cmd_mux_002|src_payload~17_combout ),
	.src_payload18(\mm_interconnect_0|cmd_mux_002|src_payload~18_combout ),
	.src_payload19(\mm_interconnect_0|cmd_mux_002|src_payload~19_combout ),
	.src_payload20(\mm_interconnect_0|cmd_mux_002|src_payload~20_combout ),
	.src_payload21(\mm_interconnect_0|cmd_mux_002|src_payload~21_combout ),
	.src_payload22(\mm_interconnect_0|cmd_mux_002|src_payload~22_combout ),
	.src_payload23(\mm_interconnect_0|cmd_mux_002|src_payload~23_combout ),
	.src_payload24(\mm_interconnect_0|cmd_mux_002|src_payload~24_combout ),
	.src_payload25(\mm_interconnect_0|cmd_mux_002|src_payload~25_combout ),
	.src_payload26(\mm_interconnect_0|cmd_mux_002|src_payload~26_combout ),
	.src_payload27(\mm_interconnect_0|cmd_mux_002|src_payload~27_combout ),
	.src_payload28(\mm_interconnect_0|cmd_mux_002|src_payload~28_combout ),
	.src_payload29(\mm_interconnect_0|cmd_mux_002|src_payload~29_combout ),
	.src_payload30(\mm_interconnect_0|cmd_mux_002|src_payload~30_combout ),
	.src_payload31(\mm_interconnect_0|cmd_mux_002|src_payload~31_combout ),
	.clk_clk(\clk_clk~input_o ));

embedded_system_altera_reset_controller rst_controller(
	.r_sync_rst1(\rst_controller|r_sync_rst~q ),
	.r_early_rst1(\rst_controller|r_early_rst~q ),
	.resetrequest(\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_oci_debug|resetrequest~q ),
	.altera_reset_synchronizer_int_chain_1(\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.clk_clk(\clk_clk~input_o ));

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 64'hEDDEFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .lut_mask = 64'hEFFFFFEFEFFFFFEF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .lut_mask = 64'hFFFFFFF7FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~0 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~1_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .lut_mask = 64'hFFFFFFFF7FFFF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[1][0]~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~3 .shared_arith = "off";

assign \clk_clk~input_o  = clk_clk;

assign ad9833_io_readdata[0] = \ad9833_comp_0|aif|good_to_reset_go~q ;

assign ad9833_io_readdata[1] = \ad9833_comp_0|aif|send_complete~q ;

assign ad9833_io_readdata[2] = \ad9833_comp_0|aif|fsync~q ;

assign ad9833_io_readdata[3] = \ad9833_comp_0|aif|sclk~q ;

assign ad9833_io_readdata[4] = \ad9833_comp_0|aif|sdata~q ;

assign ad9833_io_readdata[5] = gnd;

assign ad9833_io_readdata[6] = gnd;

assign ad9833_io_readdata[7] = gnd;

assign ad9833_io_readdata[8] = gnd;

assign ad9833_io_readdata[9] = gnd;

assign ad9833_io_readdata[10] = gnd;

assign ad9833_io_readdata[11] = gnd;

assign ad9833_io_readdata[12] = gnd;

assign ad9833_io_readdata[13] = gnd;

assign ad9833_io_readdata[14] = gnd;

assign ad9833_io_readdata[15] = gnd;

assign ad9833_io_readdata[16] = gnd;

assign ad9833_io_readdata[17] = gnd;

assign ad9833_io_readdata[18] = gnd;

assign ad9833_io_readdata[19] = gnd;

assign ad9833_io_readdata[20] = gnd;

assign ad9833_io_readdata[21] = gnd;

assign ad9833_io_readdata[22] = gnd;

assign ad9833_io_readdata[23] = gnd;

assign ad9833_io_readdata[24] = gnd;

assign ad9833_io_readdata[25] = gnd;

assign ad9833_io_readdata[26] = gnd;

assign ad9833_io_readdata[27] = gnd;

assign ad9833_io_readdata[28] = gnd;

assign ad9833_io_readdata[29] = gnd;

assign ad9833_io_readdata[30] = gnd;

assign ad9833_io_readdata[31] = gnd;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cyclonev_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 64'h6666666666666666;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 64'h9696969696969696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 64'hFFFFFFEFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 (
	.dataa(!\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\rst_controller|alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain[1]~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.dataf(!\altera_internal_jtag~TDIUTAP ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .lut_mask = 64'hEFFEFAFCEFFEFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BWHK8171:14:QXXQ6833_1~combout ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 (
	.clk(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .lut_mask = 64'h6666666666666666;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .lut_mask = 64'h6666666666666666;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .lut_mask = 64'h9696969696969696;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datac(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .lut_mask = 64'h6996966996696996;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .lut_mask = 64'h5555555555555555;
defparam \nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~4 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5 .lut_mask = 64'hFFFFFFFF7FFFF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~4 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .lut_mask = 64'hFFFFEFFFFFFFFFEF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~14_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6 .lut_mask = 64'hFFF7FFFFFFF7FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][0]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_irf_reg[2][1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~6_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .lut_mask = 64'hDEDEDEDEDEDEDEDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .lut_mask = 64'hEDDEEDDEEDDEEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .lut_mask = 64'hDEEDEDDEDEEDEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .lut_mask = 64'hEDDEDEEDDEEDEDDE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .lut_mask = 64'hBEEBEBBEBEEBEBBE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.datad(!\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_1 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_2 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\altera_internal_jtag~TDIUTAP ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 64'hFFFFB77BFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 64'hFFFFFFDFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|AMGP4450~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|AMGP4450 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|NJQG9082~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|NJQG9082 (
	.clk(\nabboc|pzdyqx_impl_inst|stratixiii_BITP7563_gen_0:stratixiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datae(!\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~4_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .lut_mask = 64'hFFFFFFDFFFFFFFDF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(!\altera_internal_jtag~TMSUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .lut_mask = 64'hFFFFFFACFFFFFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .lut_mask = 64'hDF1FDF1FDF1FDF1F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 64'hFDDFFFFFDFFDFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 64'hCF5FFFFFCF5FFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datae(!\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|ir_out[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~2_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .lut_mask = 64'hFF3F7F7FFF3F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .lut_mask = 64'hBBBBEEEEBBBBEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .lut_mask = 64'hFFFFFFFFBEEBEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .lut_mask = 64'hFFFFFFFFFFEFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(gnd),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .lut_mask = 64'hEBEBBEBEEBEBBEBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 64'h6996699669966996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .lut_mask = 64'hF7D5FFFFF7D5FFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~5 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 64'hFFFFD8FFFFFFD8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .extended_lut = "on";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .lut_mask = 64'hFF7FFFF7FF7FFFF7;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .lut_mask = 64'hFF96FF96FF96FF96;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~2_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~5_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .lut_mask = 64'h7777777777777777;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~5_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3 .lut_mask = 64'hFFFF7FF7FFFF7FF7;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2 .lut_mask = 64'h6996699669966996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~1 .lut_mask = 64'h9669699696696996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~1 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~1_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .lut_mask = 64'hFFFFFFF7FFFFFFF7;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~1 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~1 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~1 .lut_mask = 64'hFF7BFF7BFF7BFF7B;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~1 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~2 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~2 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~2 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(!\altera_internal_jtag~TDIUTAP ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .lut_mask = 64'hFBFEFBFEFBFEFBFE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .shared_arith = "off";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|comb~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|comb~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|comb~0 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \nabboc|pzdyqx_impl_inst|comb~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~0_combout ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~1_combout ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~2_combout ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .lut_mask = 64'hFBFEBFEFFBFEBFEF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 (
	.dataa(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datag(!\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .extended_lut = "on";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .lut_mask = 64'h9F6FF9F69F6FF9F6;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~12_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|Equal0~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[2][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datae(!\altera_internal_jtag~TDIUTAP ),
	.dataf(!\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .lut_mask = 64'hB1FFFFFFFFFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0 .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|sdr (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|sdr .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|sdr .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \nabboc|pzdyqx_impl_inst|sdr .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.asdata(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\nabboc|pzdyqx_impl_inst|sdr~combout ),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|dr_scan (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_1[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|dr_scan .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|dr_scan .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \nabboc|pzdyqx_impl_inst|dr_scan .shared_arith = "off";

dffeas \nabboc|pzdyqx_impl_inst|KNOR6738 (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .power_up = "low";

cyclonev_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~0 (
	.dataa(!\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.datab(!\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.datac(!\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datad(!\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.datae(!\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .extended_lut = "off";
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datad(!\nios2_qsys_0|the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[0]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_tdo_sel_reg[1]~q ),
	.dataf(!\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 64'h4747474747474747;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 64'h7777777777777777;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .lut_mask = 64'hAAAAAAAAFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .lut_mask = 64'h66666666FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(gnd),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .lut_mask = 64'h99669966FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(gnd),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .lut_mask = 64'h66999966FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .lut_mask = 64'h96696996FFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 64'h9669699696696996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 64'h7BB7B77B7BB7B77B;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal11~0_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .lut_mask = 64'h7BB7B77B7BB7B77B;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(!\altera_internal_jtag~TDIUTAP ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~3_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .lut_mask = 64'h2727272727272727;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[6]~q ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~3_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~4_combout ),
	.dataf(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .lut_mask = 64'hFFFFFFFFFFFBFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6 .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.datab(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~0_combout ),
	.datac(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~1_combout ),
	.datad(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~2_combout ),
	.datae(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7 .shared_arith = "off";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_mux_out~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cyclonev_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|~GND~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|~GND .extended_lut = "off";
defparam \auto_hub|~GND .lut_mask = 64'h0000000000000000;
defparam \auto_hub|~GND .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .shared_arith = "off";

cyclonev_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .extended_lut = "off";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:with_jtag_input_gen:instrumentation_fabric|instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .shared_arith = "off";

endmodule

module embedded_system_ad9833_avalon (
	fsync,
	good_to_reset_go,
	send_complete,
	sclk,
	sdata,
	r_sync_rst,
	wait_latency_counter_1,
	wait_latency_counter_0,
	m0_write,
	d_writedata_11,
	d_byteenable_0,
	d_writedata_10,
	d_writedata_9,
	d_writedata_8,
	d_writedata_13,
	d_writedata_12,
	d_writedata_21,
	d_writedata_20,
	d_writedata_25,
	d_writedata_17,
	d_writedata_24,
	d_writedata_16,
	d_writedata_27,
	d_writedata_19,
	d_writedata_26,
	d_writedata_18,
	d_writedata_23,
	d_writedata_15,
	d_writedata_22,
	d_writedata_14,
	d_byteenable_1,
	d_writedata_2,
	d_writedata_0,
	d_writedata_3,
	d_writedata_1,
	d_writedata_6,
	d_writedata_4,
	d_writedata_7,
	d_writedata_5,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	fsync;
output 	good_to_reset_go;
output 	send_complete;
output 	sclk;
output 	sdata;
input 	r_sync_rst;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	m0_write;
input 	d_writedata_11;
input 	d_byteenable_0;
input 	d_writedata_10;
input 	d_writedata_9;
input 	d_writedata_8;
input 	d_writedata_13;
input 	d_writedata_12;
input 	d_writedata_21;
input 	d_writedata_20;
input 	d_writedata_25;
input 	d_writedata_17;
input 	d_writedata_24;
input 	d_writedata_16;
input 	d_writedata_27;
input 	d_writedata_19;
input 	d_writedata_26;
input 	d_writedata_18;
input 	d_writedata_23;
input 	d_writedata_15;
input 	d_writedata_22;
input 	d_writedata_14;
input 	d_byteenable_1;
input 	d_writedata_2;
input 	d_writedata_0;
input 	d_writedata_3;
input 	d_writedata_1;
input 	d_writedata_6;
input 	d_writedata_4;
input 	d_writedata_7;
input 	d_writedata_5;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_ad9833if aif(
	.fsync1(fsync),
	.good_to_reset_go1(good_to_reset_go),
	.send_complete1(send_complete),
	.sclk1(sclk),
	.sdata1(sdata),
	.resetn(r_sync_rst),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.m0_write(m0_write),
	.d_writedata_11(d_writedata_11),
	.d_byteenable_0(d_byteenable_0),
	.d_writedata_10(d_writedata_10),
	.d_writedata_9(d_writedata_9),
	.d_writedata_8(d_writedata_8),
	.d_writedata_13(d_writedata_13),
	.d_writedata_12(d_writedata_12),
	.d_writedata_21(d_writedata_21),
	.d_writedata_20(d_writedata_20),
	.d_writedata_25(d_writedata_25),
	.d_writedata_17(d_writedata_17),
	.d_writedata_24(d_writedata_24),
	.d_writedata_16(d_writedata_16),
	.d_writedata_27(d_writedata_27),
	.d_writedata_19(d_writedata_19),
	.d_writedata_26(d_writedata_26),
	.d_writedata_18(d_writedata_18),
	.d_writedata_23(d_writedata_23),
	.d_writedata_15(d_writedata_15),
	.d_writedata_22(d_writedata_22),
	.d_writedata_14(d_writedata_14),
	.d_byteenable_1(d_byteenable_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_0(d_writedata_0),
	.d_writedata_3(d_writedata_3),
	.d_writedata_1(d_writedata_1),
	.d_writedata_6(d_writedata_6),
	.d_writedata_4(d_writedata_4),
	.d_writedata_7(d_writedata_7),
	.d_writedata_5(d_writedata_5),
	.clk(clk_clk));

endmodule

module embedded_system_ad9833if (
	fsync1,
	good_to_reset_go1,
	send_complete1,
	sclk1,
	sdata1,
	resetn,
	wait_latency_counter_1,
	wait_latency_counter_0,
	m0_write,
	d_writedata_11,
	d_byteenable_0,
	d_writedata_10,
	d_writedata_9,
	d_writedata_8,
	d_writedata_13,
	d_writedata_12,
	d_writedata_21,
	d_writedata_20,
	d_writedata_25,
	d_writedata_17,
	d_writedata_24,
	d_writedata_16,
	d_writedata_27,
	d_writedata_19,
	d_writedata_26,
	d_writedata_18,
	d_writedata_23,
	d_writedata_15,
	d_writedata_22,
	d_writedata_14,
	d_byteenable_1,
	d_writedata_2,
	d_writedata_0,
	d_writedata_3,
	d_writedata_1,
	d_writedata_6,
	d_writedata_4,
	d_writedata_7,
	d_writedata_5,
	clk)/* synthesis synthesis_greybox=1 */;
output 	fsync1;
output 	good_to_reset_go1;
output 	send_complete1;
output 	sclk1;
output 	sdata1;
input 	resetn;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	m0_write;
input 	d_writedata_11;
input 	d_byteenable_0;
input 	d_writedata_10;
input 	d_writedata_9;
input 	d_writedata_8;
input 	d_writedata_13;
input 	d_writedata_12;
input 	d_writedata_21;
input 	d_writedata_20;
input 	d_writedata_25;
input 	d_writedata_17;
input 	d_writedata_24;
input 	d_writedata_16;
input 	d_writedata_27;
input 	d_writedata_19;
input 	d_writedata_26;
input 	d_writedata_18;
input 	d_writedata_23;
input 	d_writedata_15;
input 	d_writedata_22;
input 	d_writedata_14;
input 	d_byteenable_1;
input 	d_writedata_2;
input 	d_writedata_0;
input 	d_writedata_3;
input 	d_writedata_1;
input 	d_writedata_6;
input 	d_writedata_4;
input 	d_writedata_7;
input 	d_writedata_5;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~25_sumout ;
wire \Add0~2 ;
wire \Add0~21_sumout ;
wire \current_node~39_combout ;
wire \current_node.0000~q ;
wire \clk_ctr[11]~2_combout ;
wire \clk_ctr[6]~q ;
wire \Add0~22 ;
wire \Add0~29_sumout ;
wire \clk_ctr[7]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \clk_ctr[8]~q ;
wire \Add0~34 ;
wire \Add0~61_sumout ;
wire \clk_ctr[9]~q ;
wire \Add0~62 ;
wire \Add0~57_sumout ;
wire \clk_ctr[10]~q ;
wire \Add0~58 ;
wire \Add0~45_sumout ;
wire \clk_ctr[11]~q ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \clk_ctr[12]~q ;
wire \Add0~50 ;
wire \Add0~37_sumout ;
wire \clk_ctr[13]~q ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \clk_ctr[14]~q ;
wire \Add0~42 ;
wire \Add0~53_sumout ;
wire \clk_ctr[15]~q ;
wire \Equal0~0_combout ;
wire \LessThan0~0_combout ;
wire \LessThan0~1_combout ;
wire \current_node~27_combout ;
wire \current_node~29_combout ;
wire \current_node~30_combout ;
wire \current_node.START_SCLK~q ;
wire \LessThan2~0_combout ;
wire \LessThan2~1_combout ;
wire \LessThan3~0_combout ;
wire \LessThan3~1_combout ;
wire \Selector28~0_combout ;
wire \Selector32~0_combout ;
wire \Selector32~1_combout ;
wire \bit_ctr[0]~q ;
wire \Selector31~0_combout ;
wire \bit_ctr[1]~q ;
wire \Selector30~0_combout ;
wire \bit_ctr[2]~q ;
wire \always0~2_combout ;
wire \Selector29~0_combout ;
wire \bit_ctr[3]~q ;
wire \always0~0_combout ;
wire \Selector28~1_combout ;
wire \bit_ctr[4]~q ;
wire \Selector27~0_combout ;
wire \bit_ctr[5]~q ;
wire \always0~1_combout ;
wire \clk_ctr[14]~0_combout ;
wire \current_node~31_combout ;
wire \Selector35~0_combout ;
wire \word_ctr[0]~q ;
wire \Selector34~0_combout ;
wire \word_ctr[1]~q ;
wire \Selector33~0_combout ;
wire \word_ctr[2]~q ;
wire \current_node~35_combout ;
wire \current_node~36_combout ;
wire \current_node.FSYNC_WAIT_LOW_1~q ;
wire \Selector2~0_combout ;
wire \current_node.START_FSYNC~q ;
wire \current_node~37_combout ;
wire \current_node~38_combout ;
wire \current_node.WORD_TRANSFER_1~q ;
wire \current_node~26_combout ;
wire \current_node~34_combout ;
wire \current_node.FSYNC_WAIT_HIGH_1~q ;
wire \current_node~32_combout ;
wire \current_node~33_combout ;
wire \current_node.SEND_COMPLETE~q ;
wire \current_node~28_combout ;
wire \current_node.CLEANUP~q ;
wire \clk_ctr[14]~1_combout ;
wire \clk_ctr[0]~q ;
wire \Add0~26 ;
wire \Add0~9_sumout ;
wire \clk_ctr[1]~q ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \clk_ctr[2]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \clk_ctr[3]~q ;
wire \Add0~18 ;
wire \Add0~5_sumout ;
wire \clk_ctr[4]~q ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \clk_ctr[5]~q ;
wire \Equal0~1_combout ;
wire \Equal0~2_combout ;
wire \Selector26~0_combout ;
wire \Selector9~0_combout ;
wire \Selector36~0_combout ;
wire \Equal4~0_combout ;
wire \Selector8~0_combout ;
wire \Equal0~3_combout ;
wire \Selector8~1_combout ;
wire \Selector8~2_combout ;
wire \Selector8~3_combout ;
wire \local_control[0]~0_combout ;
wire \local_control[10]~q ;
wire \local_control[8]~q ;
wire \local_control[9]~q ;
wire \local_control[14]~q ;
wire \local_control[12]~q ;
wire \local_control[13]~q ;
wire \local_control[15]~q ;
wire \Mux0~15_combout ;
wire \local_control[11]~q ;
wire \Mux0~0_combout ;
wire \local_freq[12]~0_combout ;
wire \local_freq[11]~q ;
wire \local_freq[10]~q ;
wire \local_freq[9]~q ;
wire \local_freq[8]~q ;
wire \Mux0~4_combout ;
wire \local_freq[13]~q ;
wire \local_freq[12]~q ;
wire \Mux0~5_combout ;
wire \local_control[2]~q ;
wire \local_control[0]~q ;
wire \local_control[1]~q ;
wire \local_control[6]~q ;
wire \local_control[4]~q ;
wire \local_control[5]~q ;
wire \local_control[7]~q ;
wire \Mux0~19_combout ;
wire \local_control[3]~q ;
wire \Mux0~6_combout ;
wire \local_freq[2]~q ;
wire \local_freq[0]~q ;
wire \local_freq[1]~q ;
wire \local_freq[6]~q ;
wire \local_freq[4]~q ;
wire \local_freq[5]~q ;
wire \local_freq[7]~q ;
wire \Mux0~23_combout ;
wire \local_freq[3]~q ;
wire \Mux0~10_combout ;
wire \Mux0~14_combout ;
wire \local_freq[21]~q ;
wire \local_freq[20]~q ;
wire \Mux2~0_combout ;
wire \local_freq[25]~q ;
wire \local_freq[17]~q ;
wire \local_freq[24]~q ;
wire \local_freq[16]~q ;
wire \Mux2~1_combout ;
wire \local_freq[27]~q ;
wire \local_freq[19]~q ;
wire \local_freq[26]~q ;
wire \local_freq[18]~q ;
wire \Mux2~2_combout ;
wire \local_freq[23]~q ;
wire \local_freq[15]~q ;
wire \local_freq[22]~q ;
wire \local_freq[14]~q ;
wire \Mux2~3_combout ;
wire \Mux2~4_combout ;
wire \sdata~0_combout ;
wire \sdata~1_combout ;


dffeas fsync(
	.clk(clk),
	.d(\Selector26~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(resetn),
	.ena(vcc),
	.q(fsync1),
	.prn(vcc));
defparam fsync.is_wysiwyg = "true";
defparam fsync.power_up = "low";

dffeas good_to_reset_go(
	.clk(clk),
	.d(\Selector9~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(good_to_reset_go1),
	.prn(vcc));
defparam good_to_reset_go.is_wysiwyg = "true";
defparam good_to_reset_go.power_up = "low";

dffeas send_complete(
	.clk(clk),
	.d(\Selector36~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(send_complete1),
	.prn(vcc));
defparam send_complete.is_wysiwyg = "true";
defparam send_complete.power_up = "low";

dffeas sclk(
	.clk(clk),
	.d(\Selector8~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(sclk1),
	.prn(vcc));
defparam sclk.is_wysiwyg = "true";
defparam sclk.power_up = "low";

dffeas sdata(
	.clk(clk),
	.d(\sdata~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sdata1),
	.prn(vcc));
defparam sdata.is_wysiwyg = "true";
defparam sdata.power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \current_node~39 (
	.dataa(!\current_node.CLEANUP~q ),
	.datab(!\current_node.0000~q ),
	.datac(!wait_latency_counter_1),
	.datad(!wait_latency_counter_0),
	.datae(!m0_write),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~39 .extended_lut = "off";
defparam \current_node~39 .lut_mask = 64'hFFFFBFFFFFFFBFFF;
defparam \current_node~39 .shared_arith = "off";

dffeas \current_node.0000 (
	.clk(clk),
	.d(\current_node~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(resetn),
	.sload(gnd),
	.ena(vcc),
	.q(\current_node.0000~q ),
	.prn(vcc));
defparam \current_node.0000 .is_wysiwyg = "true";
defparam \current_node.0000 .power_up = "low";

cyclonev_lcell_comb \clk_ctr[11]~2 (
	.dataa(!\current_node.0000~q ),
	.datab(!\current_node~28_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\clk_ctr[11]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \clk_ctr[11]~2 .extended_lut = "off";
defparam \clk_ctr[11]~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \clk_ctr[11]~2 .shared_arith = "off";

dffeas \clk_ctr[6] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[6]~q ),
	.prn(vcc));
defparam \clk_ctr[6] .is_wysiwyg = "true";
defparam \clk_ctr[6] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \clk_ctr[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[7]~q ),
	.prn(vcc));
defparam \clk_ctr[7] .is_wysiwyg = "true";
defparam \clk_ctr[7] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \clk_ctr[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[8]~q ),
	.prn(vcc));
defparam \clk_ctr[8] .is_wysiwyg = "true";
defparam \clk_ctr[8] .power_up = "low";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

dffeas \clk_ctr[9] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[9]~q ),
	.prn(vcc));
defparam \clk_ctr[9] .is_wysiwyg = "true";
defparam \clk_ctr[9] .power_up = "low";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

dffeas \clk_ctr[10] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[10]~q ),
	.prn(vcc));
defparam \clk_ctr[10] .is_wysiwyg = "true";
defparam \clk_ctr[10] .power_up = "low";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \clk_ctr[11] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[11]~q ),
	.prn(vcc));
defparam \clk_ctr[11] .is_wysiwyg = "true";
defparam \clk_ctr[11] .power_up = "low";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

dffeas \clk_ctr[12] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[12]~q ),
	.prn(vcc));
defparam \clk_ctr[12] .is_wysiwyg = "true";
defparam \clk_ctr[12] .power_up = "low";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \clk_ctr[13] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[13]~q ),
	.prn(vcc));
defparam \clk_ctr[13] .is_wysiwyg = "true";
defparam \clk_ctr[13] .power_up = "low";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \clk_ctr[14] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[14]~q ),
	.prn(vcc));
defparam \clk_ctr[14] .is_wysiwyg = "true";
defparam \clk_ctr[14] .power_up = "low";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

dffeas \clk_ctr[15] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[15]~q ),
	.prn(vcc));
defparam \clk_ctr[15] .is_wysiwyg = "true";
defparam \clk_ctr[15] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\clk_ctr[14]~q ),
	.datab(!\clk_ctr[11]~q ),
	.datac(!\clk_ctr[12]~q ),
	.datad(!\clk_ctr[15]~q ),
	.datae(!\clk_ctr[10]~q ),
	.dataf(!\clk_ctr[9]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~0 (
	.dataa(!\clk_ctr[5]~q ),
	.datab(!\clk_ctr[4]~q ),
	.datac(!\clk_ctr[6]~q ),
	.datad(!\clk_ctr[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~0 .extended_lut = "off";
defparam \LessThan0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \LessThan0~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan0~1 (
	.dataa(!\clk_ctr[8]~q ),
	.datab(!\clk_ctr[13]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\clk_ctr[2]~q ),
	.datae(!\clk_ctr[3]~q ),
	.dataf(!\LessThan0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan0~1 .extended_lut = "off";
defparam \LessThan0~1 .lut_mask = 64'hFFFFFFFFFFFFFFEF;
defparam \LessThan0~1 .shared_arith = "off";

cyclonev_lcell_comb \current_node~27 (
	.dataa(!\current_node.0000~q ),
	.datab(!wait_latency_counter_1),
	.datac(!wait_latency_counter_0),
	.datad(!m0_write),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~27 .extended_lut = "off";
defparam \current_node~27 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \current_node~27 .shared_arith = "off";

cyclonev_lcell_comb \current_node~29 (
	.dataa(!\current_node.CLEANUP~q ),
	.datab(!\current_node~28_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~29 .extended_lut = "off";
defparam \current_node~29 .lut_mask = 64'h7777777777777777;
defparam \current_node~29 .shared_arith = "off";

cyclonev_lcell_comb \current_node~30 (
	.dataa(!\current_node.START_SCLK~q ),
	.datab(!\current_node~26_combout ),
	.datac(!\LessThan0~1_combout ),
	.datad(!\current_node~27_combout ),
	.datae(!\current_node~29_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~30 .extended_lut = "off";
defparam \current_node~30 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \current_node~30 .shared_arith = "off";

dffeas \current_node.START_SCLK (
	.clk(clk),
	.d(\current_node~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_node.START_SCLK~q ),
	.prn(vcc));
defparam \current_node.START_SCLK .is_wysiwyg = "true";
defparam \current_node.START_SCLK .power_up = "low";

cyclonev_lcell_comb \LessThan2~0 (
	.dataa(!\clk_ctr[5]~q ),
	.datab(!\clk_ctr[4]~q ),
	.datac(!\clk_ctr[1]~q ),
	.datad(!\clk_ctr[0]~q ),
	.datae(!\clk_ctr[2]~q ),
	.dataf(!\clk_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~0 .extended_lut = "off";
defparam \LessThan2~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \LessThan2~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan2~1 (
	.dataa(!\clk_ctr[6]~q ),
	.datab(!\clk_ctr[7]~q ),
	.datac(!\clk_ctr[8]~q ),
	.datad(!\clk_ctr[13]~q ),
	.datae(!\Equal0~0_combout ),
	.dataf(!\LessThan2~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan2~1 .extended_lut = "off";
defparam \LessThan2~1 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \LessThan2~1 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~0 (
	.dataa(!\clk_ctr[1]~q ),
	.datab(!\clk_ctr[2]~q ),
	.datac(!\clk_ctr[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~0 .extended_lut = "off";
defparam \LessThan3~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \LessThan3~0 .shared_arith = "off";

cyclonev_lcell_comb \LessThan3~1 (
	.dataa(!\clk_ctr[8]~q ),
	.datab(!\clk_ctr[13]~q ),
	.datac(!\Equal0~0_combout ),
	.datad(!\LessThan0~0_combout ),
	.datae(!\LessThan3~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\LessThan3~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \LessThan3~1 .extended_lut = "off";
defparam \LessThan3~1 .lut_mask = 64'hFFFFFFEFFFFFFFEF;
defparam \LessThan3~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~0 (
	.dataa(!\current_node.CLEANUP~q ),
	.datab(!\current_node.WORD_TRANSFER_1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~0 .extended_lut = "off";
defparam \Selector28~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Selector28~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector32~0 (
	.dataa(!\current_node.WORD_TRANSFER_1~q ),
	.datab(!\LessThan2~1_combout ),
	.datac(!\always0~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector32~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector32~0 .extended_lut = "off";
defparam \Selector32~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector32~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector32~1 (
	.dataa(!\bit_ctr[0]~q ),
	.datab(!\LessThan3~1_combout ),
	.datac(!\Selector28~0_combout ),
	.datad(!\Selector32~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector32~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector32~1 .extended_lut = "off";
defparam \Selector32~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \Selector32~1 .shared_arith = "off";

dffeas \bit_ctr[0] (
	.clk(clk),
	.d(\Selector32~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(\bit_ctr[0]~q ),
	.prn(vcc));
defparam \bit_ctr[0] .is_wysiwyg = "true";
defparam \bit_ctr[0] .power_up = "low";

cyclonev_lcell_comb \Selector31~0 (
	.dataa(!\bit_ctr[1]~q ),
	.datab(!\bit_ctr[0]~q ),
	.datac(!\LessThan3~1_combout ),
	.datad(!\Selector28~0_combout ),
	.datae(!\Selector32~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector31~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector31~0 .extended_lut = "off";
defparam \Selector31~0 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \Selector31~0 .shared_arith = "off";

dffeas \bit_ctr[1] (
	.clk(clk),
	.d(\Selector31~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(\bit_ctr[1]~q ),
	.prn(vcc));
defparam \bit_ctr[1] .is_wysiwyg = "true";
defparam \bit_ctr[1] .power_up = "low";

cyclonev_lcell_comb \Selector30~0 (
	.dataa(!\bit_ctr[2]~q ),
	.datab(!\bit_ctr[1]~q ),
	.datac(!\bit_ctr[0]~q ),
	.datad(!\LessThan3~1_combout ),
	.datae(!\Selector28~0_combout ),
	.dataf(!\Selector32~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector30~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector30~0 .extended_lut = "off";
defparam \Selector30~0 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \Selector30~0 .shared_arith = "off";

dffeas \bit_ctr[2] (
	.clk(clk),
	.d(\Selector30~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(\bit_ctr[2]~q ),
	.prn(vcc));
defparam \bit_ctr[2] .is_wysiwyg = "true";
defparam \bit_ctr[2] .power_up = "low";

cyclonev_lcell_comb \always0~2 (
	.dataa(!\bit_ctr[2]~q ),
	.datab(!\bit_ctr[1]~q ),
	.datac(!\bit_ctr[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~2 .extended_lut = "off";
defparam \always0~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \always0~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector29~0 (
	.dataa(!\bit_ctr[3]~q ),
	.datab(!\LessThan3~1_combout ),
	.datac(!\always0~2_combout ),
	.datad(!\Selector28~0_combout ),
	.datae(!\Selector32~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector29~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector29~0 .extended_lut = "off";
defparam \Selector29~0 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \Selector29~0 .shared_arith = "off";

dffeas \bit_ctr[3] (
	.clk(clk),
	.d(\Selector29~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(\bit_ctr[3]~q ),
	.prn(vcc));
defparam \bit_ctr[3] .is_wysiwyg = "true";
defparam \bit_ctr[3] .power_up = "low";

cyclonev_lcell_comb \always0~0 (
	.dataa(!\bit_ctr[2]~q ),
	.datab(!\bit_ctr[1]~q ),
	.datac(!\bit_ctr[0]~q ),
	.datad(!\bit_ctr[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \always0~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector28~1 (
	.dataa(!\LessThan3~1_combout ),
	.datab(!\bit_ctr[4]~q ),
	.datac(!\always0~0_combout ),
	.datad(!\Selector28~0_combout ),
	.datae(!\Selector32~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector28~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector28~1 .extended_lut = "off";
defparam \Selector28~1 .lut_mask = 64'h96FFFFFF96FFFFFF;
defparam \Selector28~1 .shared_arith = "off";

dffeas \bit_ctr[4] (
	.clk(clk),
	.d(\Selector28~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(\bit_ctr[4]~q ),
	.prn(vcc));
defparam \bit_ctr[4] .is_wysiwyg = "true";
defparam \bit_ctr[4] .power_up = "low";

cyclonev_lcell_comb \Selector27~0 (
	.dataa(!\LessThan3~1_combout ),
	.datab(!\bit_ctr[5]~q ),
	.datac(!\bit_ctr[4]~q ),
	.datad(!\always0~0_combout ),
	.datae(!\Selector28~0_combout ),
	.dataf(!\Selector32~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector27~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector27~0 .extended_lut = "off";
defparam \Selector27~0 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \Selector27~0 .shared_arith = "off";

dffeas \bit_ctr[5] (
	.clk(clk),
	.d(\Selector27~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(\bit_ctr[5]~q ),
	.prn(vcc));
defparam \bit_ctr[5] .is_wysiwyg = "true";
defparam \bit_ctr[5] .power_up = "low";

cyclonev_lcell_comb \always0~1 (
	.dataa(!\bit_ctr[5]~q ),
	.datab(!\bit_ctr[4]~q ),
	.datac(!\always0~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~1 .extended_lut = "off";
defparam \always0~1 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \always0~1 .shared_arith = "off";

cyclonev_lcell_comb \clk_ctr[14]~0 (
	.dataa(!\current_node.START_SCLK~q ),
	.datab(!\current_node.FSYNC_WAIT_HIGH_1~q ),
	.datac(!\current_node.WORD_TRANSFER_1~q ),
	.datad(!\LessThan2~1_combout ),
	.datae(!\always0~1_combout ),
	.dataf(!\LessThan0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\clk_ctr[14]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \clk_ctr[14]~0 .extended_lut = "off";
defparam \clk_ctr[14]~0 .lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam \clk_ctr[14]~0 .shared_arith = "off";

cyclonev_lcell_comb \current_node~31 (
	.dataa(!\current_node.START_SCLK~q ),
	.datab(!\current_node.WORD_TRANSFER_1~q ),
	.datac(!\LessThan3~1_combout ),
	.datad(!\LessThan2~1_combout ),
	.datae(!\always0~1_combout ),
	.dataf(!\LessThan0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~31 .extended_lut = "off";
defparam \current_node~31 .lut_mask = 64'hFFFFFFFFFFFFFFF6;
defparam \current_node~31 .shared_arith = "off";

cyclonev_lcell_comb \Selector35~0 (
	.dataa(!\current_node.CLEANUP~q ),
	.datab(!\current_node.FSYNC_WAIT_LOW_1~q ),
	.datac(!\word_ctr[0]~q ),
	.datad(!\LessThan3~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector35~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector35~0 .extended_lut = "off";
defparam \Selector35~0 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \Selector35~0 .shared_arith = "off";

dffeas \word_ctr[0] (
	.clk(clk),
	.d(\Selector35~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(\word_ctr[0]~q ),
	.prn(vcc));
defparam \word_ctr[0] .is_wysiwyg = "true";
defparam \word_ctr[0] .power_up = "low";

cyclonev_lcell_comb \Selector34~0 (
	.dataa(!\current_node.CLEANUP~q ),
	.datab(!\current_node.FSYNC_WAIT_LOW_1~q ),
	.datac(!\word_ctr[0]~q ),
	.datad(!\word_ctr[1]~q ),
	.datae(!\LessThan3~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector34~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector34~0 .extended_lut = "off";
defparam \Selector34~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \Selector34~0 .shared_arith = "off";

dffeas \word_ctr[1] (
	.clk(clk),
	.d(\Selector34~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(\word_ctr[1]~q ),
	.prn(vcc));
defparam \word_ctr[1] .is_wysiwyg = "true";
defparam \word_ctr[1] .power_up = "low";

cyclonev_lcell_comb \Selector33~0 (
	.dataa(!\current_node.CLEANUP~q ),
	.datab(!\current_node.FSYNC_WAIT_LOW_1~q ),
	.datac(!\word_ctr[0]~q ),
	.datad(!\word_ctr[2]~q ),
	.datae(!\word_ctr[1]~q ),
	.dataf(!\LessThan3~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector33~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector33~0 .extended_lut = "off";
defparam \Selector33~0 .lut_mask = 64'hD77D7DD77DD7D77D;
defparam \Selector33~0 .shared_arith = "off";

dffeas \word_ctr[2] (
	.clk(clk),
	.d(\Selector33~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!resetn),
	.q(\word_ctr[2]~q ),
	.prn(vcc));
defparam \word_ctr[2] .is_wysiwyg = "true";
defparam \word_ctr[2] .power_up = "low";

cyclonev_lcell_comb \current_node~35 (
	.dataa(!\current_node.FSYNC_WAIT_HIGH_1~q ),
	.datab(!\current_node.FSYNC_WAIT_LOW_1~q ),
	.datac(!\word_ctr[2]~q ),
	.datad(!\word_ctr[1]~q ),
	.datae(!\LessThan0~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~35 .extended_lut = "off";
defparam \current_node~35 .lut_mask = 64'hFFF7FFFBFFF7FFFB;
defparam \current_node~35 .shared_arith = "off";

cyclonev_lcell_comb \current_node~36 (
	.dataa(!\current_node.FSYNC_WAIT_HIGH_1~q ),
	.datab(!\current_node.0000~q ),
	.datac(!\current_node~27_combout ),
	.datad(!\current_node~29_combout ),
	.datae(!\current_node~31_combout ),
	.dataf(!\current_node~35_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~36 .extended_lut = "off";
defparam \current_node~36 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \current_node~36 .shared_arith = "off";

dffeas \current_node.FSYNC_WAIT_LOW_1 (
	.clk(clk),
	.d(\current_node~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_node.FSYNC_WAIT_LOW_1~q ),
	.prn(vcc));
defparam \current_node.FSYNC_WAIT_LOW_1 .is_wysiwyg = "true";
defparam \current_node.FSYNC_WAIT_LOW_1 .power_up = "low";

cyclonev_lcell_comb \Selector2~0 (
	.dataa(!\current_node.START_SCLK~q ),
	.datab(!\current_node.START_FSYNC~q ),
	.datac(!\LessThan3~1_combout ),
	.datad(!\LessThan0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector2~0 .extended_lut = "off";
defparam \Selector2~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \Selector2~0 .shared_arith = "off";

dffeas \current_node.START_FSYNC (
	.clk(clk),
	.d(\Selector2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(resetn),
	.sload(gnd),
	.ena(vcc),
	.q(\current_node.START_FSYNC~q ),
	.prn(vcc));
defparam \current_node.START_FSYNC .is_wysiwyg = "true";
defparam \current_node.START_FSYNC .power_up = "low";

cyclonev_lcell_comb \current_node~37 (
	.dataa(!\current_node.FSYNC_WAIT_LOW_1~q ),
	.datab(!\current_node.START_FSYNC~q ),
	.datac(!\LessThan3~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~37 .extended_lut = "off";
defparam \current_node~37 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \current_node~37 .shared_arith = "off";

cyclonev_lcell_comb \current_node~38 (
	.dataa(!\current_node.WORD_TRANSFER_1~q ),
	.datab(!\clk_ctr[14]~0_combout ),
	.datac(!\current_node~27_combout ),
	.datad(!\current_node~29_combout ),
	.datae(!\current_node~37_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~38 .extended_lut = "off";
defparam \current_node~38 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \current_node~38 .shared_arith = "off";

dffeas \current_node.WORD_TRANSFER_1 (
	.clk(clk),
	.d(\current_node~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_node.WORD_TRANSFER_1~q ),
	.prn(vcc));
defparam \current_node.WORD_TRANSFER_1 .is_wysiwyg = "true";
defparam \current_node.WORD_TRANSFER_1 .power_up = "low";

cyclonev_lcell_comb \current_node~26 (
	.dataa(!\current_node.WORD_TRANSFER_1~q ),
	.datab(!\LessThan2~1_combout ),
	.datac(!\always0~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~26 .extended_lut = "off";
defparam \current_node~26 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \current_node~26 .shared_arith = "off";

cyclonev_lcell_comb \current_node~34 (
	.dataa(!\current_node.FSYNC_WAIT_HIGH_1~q ),
	.datab(!\current_node~26_combout ),
	.datac(!\LessThan0~1_combout ),
	.datad(!\current_node~29_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~34 .extended_lut = "off";
defparam \current_node~34 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \current_node~34 .shared_arith = "off";

dffeas \current_node.FSYNC_WAIT_HIGH_1 (
	.clk(clk),
	.d(\current_node~34_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_node.FSYNC_WAIT_HIGH_1~q ),
	.prn(vcc));
defparam \current_node.FSYNC_WAIT_HIGH_1 .is_wysiwyg = "true";
defparam \current_node.FSYNC_WAIT_HIGH_1 .power_up = "low";

cyclonev_lcell_comb \current_node~32 (
	.dataa(!\current_node.FSYNC_WAIT_HIGH_1~q ),
	.datab(!\word_ctr[2]~q ),
	.datac(!\word_ctr[1]~q ),
	.datad(!\LessThan0~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~32 .extended_lut = "off";
defparam \current_node~32 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \current_node~32 .shared_arith = "off";

cyclonev_lcell_comb \current_node~33 (
	.dataa(!\current_node.FSYNC_WAIT_HIGH_1~q ),
	.datab(!\current_node.0000~q ),
	.datac(!\current_node~27_combout ),
	.datad(!\current_node~29_combout ),
	.datae(!\current_node~31_combout ),
	.dataf(!\current_node~32_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~33 .extended_lut = "off";
defparam \current_node~33 .lut_mask = 64'hFFFFF7FFFFFFFFFF;
defparam \current_node~33 .shared_arith = "off";

dffeas \current_node.SEND_COMPLETE (
	.clk(clk),
	.d(\current_node~33_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_node.SEND_COMPLETE~q ),
	.prn(vcc));
defparam \current_node.SEND_COMPLETE .is_wysiwyg = "true";
defparam \current_node.SEND_COMPLETE .power_up = "low";

cyclonev_lcell_comb \current_node~28 (
	.dataa(!resetn),
	.datab(!\current_node.SEND_COMPLETE~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\current_node~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \current_node~28 .extended_lut = "off";
defparam \current_node~28 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \current_node~28 .shared_arith = "off";

dffeas \current_node.CLEANUP (
	.clk(clk),
	.d(\current_node~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\current_node.CLEANUP~q ),
	.prn(vcc));
defparam \current_node.CLEANUP .is_wysiwyg = "true";
defparam \current_node.CLEANUP .power_up = "low";

cyclonev_lcell_comb \clk_ctr[14]~1 (
	.dataa(!\current_node.CLEANUP~q ),
	.datab(!\current_node.FSYNC_WAIT_LOW_1~q ),
	.datac(!\current_node.START_FSYNC~q ),
	.datad(!\current_node.WORD_TRANSFER_1~q ),
	.datae(!\LessThan3~1_combout ),
	.dataf(!\clk_ctr[14]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\clk_ctr[14]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \clk_ctr[14]~1 .extended_lut = "off";
defparam \clk_ctr[14]~1 .lut_mask = 64'hFFFFBFFFFFFFFFFF;
defparam \clk_ctr[14]~1 .shared_arith = "off";

dffeas \clk_ctr[0] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[0]~q ),
	.prn(vcc));
defparam \clk_ctr[0] .is_wysiwyg = "true";
defparam \clk_ctr[0] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \clk_ctr[1] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[1]~q ),
	.prn(vcc));
defparam \clk_ctr[1] .is_wysiwyg = "true";
defparam \clk_ctr[1] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \clk_ctr[2] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[2]~q ),
	.prn(vcc));
defparam \clk_ctr[2] .is_wysiwyg = "true";
defparam \clk_ctr[2] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \clk_ctr[3] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[3]~q ),
	.prn(vcc));
defparam \clk_ctr[3] .is_wysiwyg = "true";
defparam \clk_ctr[3] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\clk_ctr[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \clk_ctr[4] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[4]~q ),
	.prn(vcc));
defparam \clk_ctr[4] .is_wysiwyg = "true";
defparam \clk_ctr[4] .power_up = "low";

dffeas \clk_ctr[5] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\clk_ctr[14]~1_combout ),
	.sload(gnd),
	.ena(\clk_ctr[11]~2_combout ),
	.q(\clk_ctr[5]~q ),
	.prn(vcc));
defparam \clk_ctr[5] .is_wysiwyg = "true";
defparam \clk_ctr[5] .power_up = "low";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!\clk_ctr[6]~q ),
	.datab(!\clk_ctr[0]~q ),
	.datac(!\clk_ctr[7]~q ),
	.datad(!\clk_ctr[8]~q ),
	.datae(!\clk_ctr[13]~q ),
	.dataf(!\Equal0~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~2 (
	.dataa(!\clk_ctr[5]~q ),
	.datab(!\clk_ctr[4]~q ),
	.datac(!\clk_ctr[1]~q ),
	.datad(!\clk_ctr[2]~q ),
	.datae(!\clk_ctr[3]~q ),
	.dataf(!\Equal0~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector26~0 (
	.dataa(!fsync1),
	.datab(!\Equal0~2_combout ),
	.datac(!\current_node.FSYNC_WAIT_HIGH_1~q ),
	.datad(!\current_node.FSYNC_WAIT_LOW_1~q ),
	.datae(!\current_node.START_FSYNC~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector26~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector26~0 .extended_lut = "off";
defparam \Selector26~0 .lut_mask = 64'hFF7FDF5FFF7FDF5F;
defparam \Selector26~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector9~0 (
	.dataa(!good_to_reset_go1),
	.datab(!\current_node.START_SCLK~q ),
	.datac(!\Equal0~2_combout ),
	.datad(!\current_node.CLEANUP~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector9~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector9~0 .extended_lut = "off";
defparam \Selector9~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \Selector9~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector36~0 (
	.dataa(!send_complete1),
	.datab(!\current_node.CLEANUP~q ),
	.datac(!\current_node.SEND_COMPLETE~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector36~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector36~0 .extended_lut = "off";
defparam \Selector36~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \Selector36~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal4~0 (
	.dataa(!\clk_ctr[5]~q ),
	.datab(!\clk_ctr[4]~q ),
	.datac(!\clk_ctr[1]~q ),
	.datad(!\clk_ctr[2]~q ),
	.datae(!\clk_ctr[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal4~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal4~0 .extended_lut = "off";
defparam \Equal4~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \Equal4~0 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~0 (
	.dataa(!\current_node.START_SCLK~q ),
	.datab(!\Equal0~1_combout ),
	.datac(!\current_node.FSYNC_WAIT_HIGH_1~q ),
	.datad(!\current_node.WORD_TRANSFER_1~q ),
	.datae(!\Equal4~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~0 .extended_lut = "off";
defparam \Selector8~0 .lut_mask = 64'hA3FFFFFFA3FFFFFF;
defparam \Selector8~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~3 (
	.dataa(!\clk_ctr[7]~q ),
	.datab(!\clk_ctr[8]~q ),
	.datac(!\clk_ctr[13]~q ),
	.datad(!\Equal0~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~3 .extended_lut = "off";
defparam \Equal0~3 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \Equal0~3 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~1 (
	.dataa(!\clk_ctr[1]~q ),
	.datab(!\clk_ctr[0]~q ),
	.datac(!\clk_ctr[2]~q ),
	.datad(!\clk_ctr[3]~q ),
	.datae(!\current_node.WORD_TRANSFER_1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~1 .extended_lut = "off";
defparam \Selector8~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \Selector8~1 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~2 (
	.dataa(!\clk_ctr[5]~q ),
	.datab(!\clk_ctr[4]~q ),
	.datac(!\clk_ctr[6]~q ),
	.datad(!\Equal0~3_combout ),
	.datae(!\Selector8~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~2 .extended_lut = "off";
defparam \Selector8~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \Selector8~2 .shared_arith = "off";

cyclonev_lcell_comb \Selector8~3 (
	.dataa(!sclk1),
	.datab(!\current_node.START_SCLK~q ),
	.datac(!\Equal0~2_combout ),
	.datad(!\current_node.WORD_TRANSFER_1~q ),
	.datae(!\Selector8~0_combout ),
	.dataf(!\Selector8~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Selector8~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Selector8~3 .extended_lut = "off";
defparam \Selector8~3 .lut_mask = 64'hF7FF37FFFFFFFFFF;
defparam \Selector8~3 .shared_arith = "off";

cyclonev_lcell_comb \local_control[0]~0 (
	.dataa(!resetn),
	.datab(!d_byteenable_0),
	.datac(!d_byteenable_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_control[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \local_control[0]~0 .extended_lut = "off";
defparam \local_control[0]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \local_control[0]~0 .shared_arith = "off";

dffeas \local_control[10] (
	.clk(clk),
	.d(d_writedata_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[10]~q ),
	.prn(vcc));
defparam \local_control[10] .is_wysiwyg = "true";
defparam \local_control[10] .power_up = "low";

dffeas \local_control[8] (
	.clk(clk),
	.d(d_writedata_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[8]~q ),
	.prn(vcc));
defparam \local_control[8] .is_wysiwyg = "true";
defparam \local_control[8] .power_up = "low";

dffeas \local_control[9] (
	.clk(clk),
	.d(d_writedata_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[9]~q ),
	.prn(vcc));
defparam \local_control[9] .is_wysiwyg = "true";
defparam \local_control[9] .power_up = "low";

dffeas \local_control[14] (
	.clk(clk),
	.d(d_writedata_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[14]~q ),
	.prn(vcc));
defparam \local_control[14] .is_wysiwyg = "true";
defparam \local_control[14] .power_up = "low";

dffeas \local_control[12] (
	.clk(clk),
	.d(d_writedata_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[12]~q ),
	.prn(vcc));
defparam \local_control[12] .is_wysiwyg = "true";
defparam \local_control[12] .power_up = "low";

dffeas \local_control[13] (
	.clk(clk),
	.d(d_writedata_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[13]~q ),
	.prn(vcc));
defparam \local_control[13] .is_wysiwyg = "true";
defparam \local_control[13] .power_up = "low";

dffeas \local_control[15] (
	.clk(clk),
	.d(d_writedata_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[15]~q ),
	.prn(vcc));
defparam \local_control[15] .is_wysiwyg = "true";
defparam \local_control[15] .power_up = "low";

cyclonev_lcell_comb \Mux0~15 (
	.dataa(!\local_control[14]~q ),
	.datab(!\local_control[12]~q ),
	.datac(!\local_control[13]~q ),
	.datad(!\bit_ctr[0]~q ),
	.datae(!\bit_ctr[1]~q ),
	.dataf(!\bit_ctr[2]~q ),
	.datag(!\local_control[15]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~15 .extended_lut = "on";
defparam \Mux0~15 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \Mux0~15 .shared_arith = "off";

dffeas \local_control[11] (
	.clk(clk),
	.d(d_writedata_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[11]~q ),
	.prn(vcc));
defparam \local_control[11] .is_wysiwyg = "true";
defparam \local_control[11] .power_up = "low";

cyclonev_lcell_comb \Mux0~0 (
	.dataa(!\local_control[10]~q ),
	.datab(!\local_control[8]~q ),
	.datac(!\local_control[9]~q ),
	.datad(!\bit_ctr[2]~q ),
	.datae(!\bit_ctr[1]~q ),
	.dataf(!\Mux0~15_combout ),
	.datag(!\local_control[11]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~0 .extended_lut = "on";
defparam \Mux0~0 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \Mux0~0 .shared_arith = "off";

cyclonev_lcell_comb \local_freq[12]~0 (
	.dataa(!resetn),
	.datab(!d_byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\local_freq[12]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \local_freq[12]~0 .extended_lut = "off";
defparam \local_freq[12]~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \local_freq[12]~0 .shared_arith = "off";

dffeas \local_freq[11] (
	.clk(clk),
	.d(d_writedata_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[11]~q ),
	.prn(vcc));
defparam \local_freq[11] .is_wysiwyg = "true";
defparam \local_freq[11] .power_up = "low";

dffeas \local_freq[10] (
	.clk(clk),
	.d(d_writedata_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[10]~q ),
	.prn(vcc));
defparam \local_freq[10] .is_wysiwyg = "true";
defparam \local_freq[10] .power_up = "low";

dffeas \local_freq[9] (
	.clk(clk),
	.d(d_writedata_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[9]~q ),
	.prn(vcc));
defparam \local_freq[9] .is_wysiwyg = "true";
defparam \local_freq[9] .power_up = "low";

dffeas \local_freq[8] (
	.clk(clk),
	.d(d_writedata_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[8]~q ),
	.prn(vcc));
defparam \local_freq[8] .is_wysiwyg = "true";
defparam \local_freq[8] .power_up = "low";

cyclonev_lcell_comb \Mux0~4 (
	.dataa(!\local_freq[11]~q ),
	.datab(!\local_freq[10]~q ),
	.datac(!\local_freq[9]~q ),
	.datad(!\local_freq[8]~q ),
	.datae(!\bit_ctr[0]~q ),
	.dataf(!\bit_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~4 .extended_lut = "off";
defparam \Mux0~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux0~4 .shared_arith = "off";

dffeas \local_freq[13] (
	.clk(clk),
	.d(d_writedata_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[13]~q ),
	.prn(vcc));
defparam \local_freq[13] .is_wysiwyg = "true";
defparam \local_freq[13] .power_up = "low";

dffeas \local_freq[12] (
	.clk(clk),
	.d(d_writedata_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[12]~q ),
	.prn(vcc));
defparam \local_freq[12] .is_wysiwyg = "true";
defparam \local_freq[12] .power_up = "low";

cyclonev_lcell_comb \Mux0~5 (
	.dataa(!\bit_ctr[2]~q ),
	.datab(!\bit_ctr[1]~q ),
	.datac(!\bit_ctr[0]~q ),
	.datad(!\Mux0~4_combout ),
	.datae(!\local_freq[13]~q ),
	.dataf(!\local_freq[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~5 .extended_lut = "off";
defparam \Mux0~5 .lut_mask = 64'h96FFFFFFFFFFFFFF;
defparam \Mux0~5 .shared_arith = "off";

dffeas \local_control[2] (
	.clk(clk),
	.d(d_writedata_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[2]~q ),
	.prn(vcc));
defparam \local_control[2] .is_wysiwyg = "true";
defparam \local_control[2] .power_up = "low";

dffeas \local_control[0] (
	.clk(clk),
	.d(d_writedata_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[0]~q ),
	.prn(vcc));
defparam \local_control[0] .is_wysiwyg = "true";
defparam \local_control[0] .power_up = "low";

dffeas \local_control[1] (
	.clk(clk),
	.d(d_writedata_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[1]~q ),
	.prn(vcc));
defparam \local_control[1] .is_wysiwyg = "true";
defparam \local_control[1] .power_up = "low";

dffeas \local_control[6] (
	.clk(clk),
	.d(d_writedata_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[6]~q ),
	.prn(vcc));
defparam \local_control[6] .is_wysiwyg = "true";
defparam \local_control[6] .power_up = "low";

dffeas \local_control[4] (
	.clk(clk),
	.d(d_writedata_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[4]~q ),
	.prn(vcc));
defparam \local_control[4] .is_wysiwyg = "true";
defparam \local_control[4] .power_up = "low";

dffeas \local_control[5] (
	.clk(clk),
	.d(d_writedata_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[5]~q ),
	.prn(vcc));
defparam \local_control[5] .is_wysiwyg = "true";
defparam \local_control[5] .power_up = "low";

dffeas \local_control[7] (
	.clk(clk),
	.d(d_writedata_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[7]~q ),
	.prn(vcc));
defparam \local_control[7] .is_wysiwyg = "true";
defparam \local_control[7] .power_up = "low";

cyclonev_lcell_comb \Mux0~19 (
	.dataa(!\local_control[6]~q ),
	.datab(!\local_control[4]~q ),
	.datac(!\local_control[5]~q ),
	.datad(!\bit_ctr[0]~q ),
	.datae(!\bit_ctr[1]~q ),
	.dataf(!\bit_ctr[2]~q ),
	.datag(!\local_control[7]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~19 .extended_lut = "on";
defparam \Mux0~19 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \Mux0~19 .shared_arith = "off";

dffeas \local_control[3] (
	.clk(clk),
	.d(d_writedata_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_control[0]~0_combout ),
	.q(\local_control[3]~q ),
	.prn(vcc));
defparam \local_control[3] .is_wysiwyg = "true";
defparam \local_control[3] .power_up = "low";

cyclonev_lcell_comb \Mux0~6 (
	.dataa(!\local_control[2]~q ),
	.datab(!\local_control[0]~q ),
	.datac(!\local_control[1]~q ),
	.datad(!\bit_ctr[2]~q ),
	.datae(!\bit_ctr[1]~q ),
	.dataf(!\Mux0~19_combout ),
	.datag(!\local_control[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~6 .extended_lut = "on";
defparam \Mux0~6 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \Mux0~6 .shared_arith = "off";

dffeas \local_freq[2] (
	.clk(clk),
	.d(d_writedata_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[2]~q ),
	.prn(vcc));
defparam \local_freq[2] .is_wysiwyg = "true";
defparam \local_freq[2] .power_up = "low";

dffeas \local_freq[0] (
	.clk(clk),
	.d(d_writedata_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[0]~q ),
	.prn(vcc));
defparam \local_freq[0] .is_wysiwyg = "true";
defparam \local_freq[0] .power_up = "low";

dffeas \local_freq[1] (
	.clk(clk),
	.d(d_writedata_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[1]~q ),
	.prn(vcc));
defparam \local_freq[1] .is_wysiwyg = "true";
defparam \local_freq[1] .power_up = "low";

dffeas \local_freq[6] (
	.clk(clk),
	.d(d_writedata_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[6]~q ),
	.prn(vcc));
defparam \local_freq[6] .is_wysiwyg = "true";
defparam \local_freq[6] .power_up = "low";

dffeas \local_freq[4] (
	.clk(clk),
	.d(d_writedata_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[4]~q ),
	.prn(vcc));
defparam \local_freq[4] .is_wysiwyg = "true";
defparam \local_freq[4] .power_up = "low";

dffeas \local_freq[5] (
	.clk(clk),
	.d(d_writedata_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[5]~q ),
	.prn(vcc));
defparam \local_freq[5] .is_wysiwyg = "true";
defparam \local_freq[5] .power_up = "low";

dffeas \local_freq[7] (
	.clk(clk),
	.d(d_writedata_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[7]~q ),
	.prn(vcc));
defparam \local_freq[7] .is_wysiwyg = "true";
defparam \local_freq[7] .power_up = "low";

cyclonev_lcell_comb \Mux0~23 (
	.dataa(!\local_freq[6]~q ),
	.datab(!\local_freq[4]~q ),
	.datac(!\local_freq[5]~q ),
	.datad(!\bit_ctr[0]~q ),
	.datae(!\bit_ctr[1]~q ),
	.dataf(!\bit_ctr[2]~q ),
	.datag(!\local_freq[7]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~23 .extended_lut = "on";
defparam \Mux0~23 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \Mux0~23 .shared_arith = "off";

dffeas \local_freq[3] (
	.clk(clk),
	.d(d_writedata_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[3]~q ),
	.prn(vcc));
defparam \local_freq[3] .is_wysiwyg = "true";
defparam \local_freq[3] .power_up = "low";

cyclonev_lcell_comb \Mux0~10 (
	.dataa(!\local_freq[2]~q ),
	.datab(!\local_freq[0]~q ),
	.datac(!\local_freq[1]~q ),
	.datad(!\bit_ctr[2]~q ),
	.datae(!\bit_ctr[1]~q ),
	.dataf(!\Mux0~23_combout ),
	.datag(!\local_freq[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~10 .extended_lut = "on";
defparam \Mux0~10 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \Mux0~10 .shared_arith = "off";

cyclonev_lcell_comb \Mux0~14 (
	.dataa(!\Mux0~0_combout ),
	.datab(!\Mux0~5_combout ),
	.datac(!\Mux0~6_combout ),
	.datad(!\Mux0~10_combout ),
	.datae(!\word_ctr[0]~q ),
	.dataf(!\bit_ctr[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux0~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux0~14 .extended_lut = "off";
defparam \Mux0~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux0~14 .shared_arith = "off";

dffeas \local_freq[21] (
	.clk(clk),
	.d(d_writedata_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[21]~q ),
	.prn(vcc));
defparam \local_freq[21] .is_wysiwyg = "true";
defparam \local_freq[21] .power_up = "low";

dffeas \local_freq[20] (
	.clk(clk),
	.d(d_writedata_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[20]~q ),
	.prn(vcc));
defparam \local_freq[20] .is_wysiwyg = "true";
defparam \local_freq[20] .power_up = "low";

cyclonev_lcell_comb \Mux2~0 (
	.dataa(!\bit_ctr[0]~q ),
	.datab(!\bit_ctr[3]~q ),
	.datac(!\local_freq[21]~q ),
	.datad(!\local_freq[20]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~0 .extended_lut = "off";
defparam \Mux2~0 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \Mux2~0 .shared_arith = "off";

dffeas \local_freq[25] (
	.clk(clk),
	.d(d_writedata_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[25]~q ),
	.prn(vcc));
defparam \local_freq[25] .is_wysiwyg = "true";
defparam \local_freq[25] .power_up = "low";

dffeas \local_freq[17] (
	.clk(clk),
	.d(d_writedata_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[17]~q ),
	.prn(vcc));
defparam \local_freq[17] .is_wysiwyg = "true";
defparam \local_freq[17] .power_up = "low";

dffeas \local_freq[24] (
	.clk(clk),
	.d(d_writedata_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[24]~q ),
	.prn(vcc));
defparam \local_freq[24] .is_wysiwyg = "true";
defparam \local_freq[24] .power_up = "low";

dffeas \local_freq[16] (
	.clk(clk),
	.d(d_writedata_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[16]~q ),
	.prn(vcc));
defparam \local_freq[16] .is_wysiwyg = "true";
defparam \local_freq[16] .power_up = "low";

cyclonev_lcell_comb \Mux2~1 (
	.dataa(!\local_freq[25]~q ),
	.datab(!\local_freq[17]~q ),
	.datac(!\local_freq[24]~q ),
	.datad(!\local_freq[16]~q ),
	.datae(!\bit_ctr[3]~q ),
	.dataf(!\bit_ctr[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~1 .extended_lut = "off";
defparam \Mux2~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~1 .shared_arith = "off";

dffeas \local_freq[27] (
	.clk(clk),
	.d(d_writedata_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[27]~q ),
	.prn(vcc));
defparam \local_freq[27] .is_wysiwyg = "true";
defparam \local_freq[27] .power_up = "low";

dffeas \local_freq[19] (
	.clk(clk),
	.d(d_writedata_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[19]~q ),
	.prn(vcc));
defparam \local_freq[19] .is_wysiwyg = "true";
defparam \local_freq[19] .power_up = "low";

dffeas \local_freq[26] (
	.clk(clk),
	.d(d_writedata_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[26]~q ),
	.prn(vcc));
defparam \local_freq[26] .is_wysiwyg = "true";
defparam \local_freq[26] .power_up = "low";

dffeas \local_freq[18] (
	.clk(clk),
	.d(d_writedata_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[18]~q ),
	.prn(vcc));
defparam \local_freq[18] .is_wysiwyg = "true";
defparam \local_freq[18] .power_up = "low";

cyclonev_lcell_comb \Mux2~2 (
	.dataa(!\local_freq[27]~q ),
	.datab(!\local_freq[19]~q ),
	.datac(!\local_freq[26]~q ),
	.datad(!\local_freq[18]~q ),
	.datae(!\bit_ctr[3]~q ),
	.dataf(!\bit_ctr[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~2 .extended_lut = "off";
defparam \Mux2~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~2 .shared_arith = "off";

dffeas \local_freq[23] (
	.clk(clk),
	.d(d_writedata_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[23]~q ),
	.prn(vcc));
defparam \local_freq[23] .is_wysiwyg = "true";
defparam \local_freq[23] .power_up = "low";

dffeas \local_freq[15] (
	.clk(clk),
	.d(d_writedata_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[15]~q ),
	.prn(vcc));
defparam \local_freq[15] .is_wysiwyg = "true";
defparam \local_freq[15] .power_up = "low";

dffeas \local_freq[22] (
	.clk(clk),
	.d(d_writedata_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[22]~q ),
	.prn(vcc));
defparam \local_freq[22] .is_wysiwyg = "true";
defparam \local_freq[22] .power_up = "low";

dffeas \local_freq[14] (
	.clk(clk),
	.d(d_writedata_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\local_freq[12]~0_combout ),
	.q(\local_freq[14]~q ),
	.prn(vcc));
defparam \local_freq[14] .is_wysiwyg = "true";
defparam \local_freq[14] .power_up = "low";

cyclonev_lcell_comb \Mux2~3 (
	.dataa(!\local_freq[23]~q ),
	.datab(!\local_freq[15]~q ),
	.datac(!\local_freq[22]~q ),
	.datad(!\local_freq[14]~q ),
	.datae(!\bit_ctr[3]~q ),
	.dataf(!\bit_ctr[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~3 .extended_lut = "off";
defparam \Mux2~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~3 .shared_arith = "off";

cyclonev_lcell_comb \Mux2~4 (
	.dataa(!\Mux2~0_combout ),
	.datab(!\Mux2~1_combout ),
	.datac(!\Mux2~2_combout ),
	.datad(!\Mux2~3_combout ),
	.datae(!\bit_ctr[2]~q ),
	.dataf(!\bit_ctr[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux2~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux2~4 .extended_lut = "off";
defparam \Mux2~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \Mux2~4 .shared_arith = "off";

cyclonev_lcell_comb \sdata~0 (
	.dataa(!\Mux0~14_combout ),
	.datab(!\word_ctr[2]~q ),
	.datac(!\word_ctr[1]~q ),
	.datad(!\Mux2~4_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdata~0 .extended_lut = "off";
defparam \sdata~0 .lut_mask = 64'h7DFF7DFF7DFF7DFF;
defparam \sdata~0 .shared_arith = "off";

cyclonev_lcell_comb \sdata~1 (
	.dataa(!sdata1),
	.datab(!\Equal0~2_combout ),
	.datac(!resetn),
	.datad(!\current_node.WORD_TRANSFER_1~q ),
	.datae(!\sdata~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sdata~1 .extended_lut = "off";
defparam \sdata~1 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \sdata~1 .shared_arith = "off";

endmodule

module embedded_system_altera_reset_controller (
	r_sync_rst1,
	r_early_rst1,
	resetrequest,
	altera_reset_synchronizer_int_chain_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	r_sync_rst1;
output 	r_early_rst1;
input 	resetrequest;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;
wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[2]~q ;
wire \altera_reset_synchronizer_int_chain[3]~q ;
wire \altera_reset_synchronizer_int_chain[4]~0_combout ;
wire \altera_reset_synchronizer_int_chain[4]~q ;
wire \r_sync_rst_chain[3]~q ;
wire \r_sync_rst_chain~1_combout ;
wire \r_sync_rst_chain[2]~q ;
wire \r_sync_rst_chain~0_combout ;
wire \r_sync_rst_chain[1]~q ;
wire \WideOr0~0_combout ;
wire \always2~0_combout ;


embedded_system_altera_reset_synchronizer alt_rst_req_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.altera_reset_synchronizer_int_chain_1(altera_reset_synchronizer_int_chain_1),
	.clk(clk_clk));

embedded_system_altera_reset_synchronizer_1 alt_rst_sync_uq1(
	.altera_reset_synchronizer_int_chain_out1(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.resetrequest(resetrequest),
	.clk(clk_clk));

dffeas r_sync_rst(
	.clk(clk_clk),
	.d(\WideOr0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_sync_rst1),
	.prn(vcc));
defparam r_sync_rst.is_wysiwyg = "true";
defparam r_sync_rst.power_up = "low";

dffeas r_early_rst(
	.clk(clk_clk),
	.d(\always2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(r_early_rst1),
	.prn(vcc));
defparam r_early_rst.is_wysiwyg = "true";
defparam r_early_rst.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk_clk),
	.d(\alt_rst_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[2] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[2]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[2] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[2] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[3]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[3] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[3] .power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[4]~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[4]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[4]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \altera_reset_synchronizer_int_chain[4]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[4] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[4]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[4]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[4] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[4] .power_up = "low";

dffeas \r_sync_rst_chain[3] (
	.clk(clk_clk),
	.d(\altera_reset_synchronizer_int_chain[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[3]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[3] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[3] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~1 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~1 .extended_lut = "off";
defparam \r_sync_rst_chain~1 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~1 .shared_arith = "off";

dffeas \r_sync_rst_chain[2] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[2]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[2] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[2] .power_up = "low";

cyclonev_lcell_comb \r_sync_rst_chain~0 (
	.dataa(!\altera_reset_synchronizer_int_chain[2]~q ),
	.datab(!\r_sync_rst_chain[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\r_sync_rst_chain~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \r_sync_rst_chain~0 .extended_lut = "off";
defparam \r_sync_rst_chain~0 .lut_mask = 64'h7777777777777777;
defparam \r_sync_rst_chain~0 .shared_arith = "off";

dffeas \r_sync_rst_chain[1] (
	.clk(clk_clk),
	.d(\r_sync_rst_chain~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\r_sync_rst_chain[1]~q ),
	.prn(vcc));
defparam \r_sync_rst_chain[1] .is_wysiwyg = "true";
defparam \r_sync_rst_chain[1] .power_up = "low";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!r_sync_rst1),
	.datab(!\altera_reset_synchronizer_int_chain[4]~q ),
	.datac(!\r_sync_rst_chain[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\WideOr0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \always2~0 (
	.dataa(!\r_sync_rst_chain[2]~q ),
	.datab(!\alt_rst_req_sync_uq1|altera_reset_synchronizer_int_chain_out~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always2~0 .extended_lut = "off";
defparam \always2~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \always2~0 .shared_arith = "off";

endmodule

module embedded_system_altera_reset_synchronizer (
	altera_reset_synchronizer_int_chain_out1,
	altera_reset_synchronizer_int_chain_1,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
output 	altera_reset_synchronizer_int_chain_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

cyclonev_lcell_comb \altera_reset_synchronizer_int_chain[1]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(altera_reset_synchronizer_int_chain_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \altera_reset_synchronizer_int_chain[1]~0 .extended_lut = "off";
defparam \altera_reset_synchronizer_int_chain[1]~0 .lut_mask = 64'h0000000000000000;
defparam \altera_reset_synchronizer_int_chain[1]~0 .shared_arith = "off";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(altera_reset_synchronizer_int_chain_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module embedded_system_altera_reset_synchronizer_1 (
	altera_reset_synchronizer_int_chain_out1,
	resetrequest,
	clk)/* synthesis synthesis_greybox=1 */;
output 	altera_reset_synchronizer_int_chain_out1;
input 	resetrequest;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \altera_reset_synchronizer_int_chain[1]~q ;
wire \altera_reset_synchronizer_int_chain[0]~q ;


dffeas altera_reset_synchronizer_int_chain_out(
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[0]~q ),
	.asdata(vcc),
	.clrn(!resetrequest),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(altera_reset_synchronizer_int_chain_out1),
	.prn(vcc));
defparam altera_reset_synchronizer_int_chain_out.is_wysiwyg = "true";
defparam altera_reset_synchronizer_int_chain_out.power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!resetrequest),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[1]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[1] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[1] .power_up = "low";

dffeas \altera_reset_synchronizer_int_chain[0] (
	.clk(clk),
	.d(\altera_reset_synchronizer_int_chain[1]~q ),
	.asdata(vcc),
	.clrn(!resetrequest),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\altera_reset_synchronizer_int_chain[0]~q ),
	.prn(vcc));
defparam \altera_reset_synchronizer_int_chain[0] .is_wysiwyg = "true";
defparam \altera_reset_synchronizer_int_chain[0] .power_up = "low";

endmodule

module embedded_system_embedded_system_mm_interconnect_0 (
	q_a_2,
	q_a_10,
	q_a_18,
	q_a_26,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_29,
	q_a_13,
	q_a_28,
	q_a_12,
	q_a_27,
	q_a_11,
	q_a_25,
	q_a_9,
	q_a_24,
	q_a_8,
	q_a_6,
	q_a_14,
	q_a_22,
	q_a_30,
	q_a_5,
	q_a_21,
	q_a_4,
	q_a_20,
	q_a_3,
	q_a_19,
	q_a_1,
	q_a_17,
	q_a_0,
	q_a_16,
	readdata_2,
	readdata_10,
	readdata_18,
	readdata_26,
	readdata_7,
	readdata_23,
	readdata_15,
	readdata_31,
	readdata_29,
	readdata_13,
	readdata_28,
	readdata_12,
	readdata_27,
	readdata_11,
	readdata_25,
	readdata_9,
	readdata_24,
	readdata_8,
	readdata_6,
	readdata_14,
	readdata_22,
	readdata_30,
	readdata_5,
	readdata_21,
	readdata_4,
	readdata_20,
	readdata_3,
	readdata_19,
	readdata_1,
	readdata_17,
	readdata_0,
	readdata_16,
	r_sync_rst,
	wait_latency_counter_1,
	wait_latency_counter_0,
	hold_waitrequest,
	d_address_offset_field_0,
	d_write,
	d_address_tag_field_2,
	d_address_tag_field_1,
	d_address_tag_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	d_address_line_field_2,
	d_address_line_field_1,
	d_address_line_field_0,
	d_address_offset_field_2,
	d_address_offset_field_1,
	m0_write,
	d_writedata_11,
	d_byteenable_0,
	d_writedata_10,
	d_writedata_9,
	d_writedata_8,
	d_writedata_13,
	d_writedata_12,
	d_writedata_21,
	d_writedata_20,
	d_writedata_25,
	d_writedata_17,
	d_writedata_24,
	d_writedata_16,
	d_writedata_27,
	d_writedata_19,
	d_writedata_26,
	d_writedata_18,
	d_writedata_23,
	d_writedata_15,
	d_writedata_22,
	d_writedata_14,
	d_read,
	suppress_change_dest_id,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	saved_grant_01,
	mem_used_11,
	WideOr0,
	av_waitrequest,
	d_byteenable_1,
	d_writedata_2,
	d_writedata_0,
	d_writedata_3,
	d_writedata_1,
	hbreak_enabled,
	i_read,
	src0_valid,
	ic_fill_tag_1,
	ic_fill_tag_0,
	ic_fill_line_6,
	Equal1,
	src0_valid1,
	src1_valid,
	saved_grant_1,
	rf_source_valid,
	src1_valid1,
	src2_valid,
	saved_grant_11,
	d_writedata_6,
	d_writedata_4,
	d_writedata_7,
	d_writedata_5,
	WideOr1,
	suppress_change_dest_id1,
	WideOr01,
	WideOr02,
	nonposted_cmd_accepted,
	ic_fill_line_5,
	src_data_46,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	ic_fill_line_1,
	src_data_42,
	ic_fill_line_0,
	src_data_41,
	ic_fill_ap_offset_2,
	src_data_40,
	ic_fill_ap_offset_1,
	src_data_39,
	ic_fill_line_4,
	src_data_45,
	ic_fill_line_3,
	src_data_44,
	ic_fill_line_2,
	src_data_43,
	src_payload1,
	src_data_32,
	src_payload2,
	src_payload3,
	WideOr11,
	src_data_2,
	src_data_10,
	src_data_18,
	src_data_26,
	src_data_7,
	src_data_23,
	src_data_15,
	src_data_31,
	src_data_29,
	src_data_13,
	src_data_28,
	src_data_12,
	src_data_27,
	src_data_11,
	src_data_25,
	src_data_9,
	src_data_24,
	src_data_8,
	src_data_6,
	src_data_14,
	src_data_22,
	src_data_30,
	src_data_5,
	src_data_21,
	src_data_4,
	src_data_20,
	src_data_3,
	src_data_19,
	src_data_1,
	src_data_17,
	src_data_0,
	src_data_16,
	src_payload4,
	src_data_51,
	src_data_33,
	src_data_110,
	src_data_47,
	src_data_210,
	src_data_281,
	src_data_311,
	src_data_271,
	src_data_291,
	src_data_301,
	src_data_01,
	src_data_231,
	src_data_261,
	src_data_221,
	src_data_241,
	src_data_251,
	src_data_161,
	src_data_151,
	src_data_131,
	src_data_141,
	src_data_121,
	src_data_111,
	src_data_81,
	src_payload5,
	src_data_381,
	src_data_391,
	src_data_401,
	src_data_411,
	src_data_421,
	src_data_431,
	src_data_441,
	src_data_451,
	src_data_461,
	src_data_471,
	src_data_321,
	src_payload6,
	src_data_331,
	src_payload7,
	d_byteenable_2,
	src_data_34,
	src_payload8,
	d_byteenable_3,
	src_data_35,
	src_data_191,
	src_payload9,
	src_payload10,
	src_payload11,
	d_writedata_31,
	src_payload12,
	d_writedata_29,
	src_payload13,
	src_payload14,
	src_data_181,
	d_writedata_28,
	src_payload15,
	src_payload16,
	src_data_171,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	d_writedata_30,
	src_payload26,
	src_payload27,
	src_payload28,
	src_data_101,
	src_payload29,
	src_payload30,
	src_data_91,
	src_payload31,
	src_payload32,
	src_payload33,
	src_payload34,
	src_payload35,
	src_payload36,
	src_data_211,
	src_data_201,
	src_data_71,
	src_data_61,
	src_payload37,
	src_data_351,
	src_payload38,
	src_payload39,
	src_data_341,
	src_payload40,
	src_payload41,
	src_payload42,
	src_payload43,
	src_payload44,
	src_payload45,
	src_payload46,
	src_payload47,
	src_payload48,
	src_payload49,
	src_payload50,
	src_payload51,
	src_payload52,
	src_payload53,
	src_data_332,
	src_payload54,
	src_payload55,
	src_payload56,
	src_payload57,
	src_payload58,
	src_payload59,
	src_payload60,
	src_payload61,
	src_payload62,
	src_payload63,
	src_payload64,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	q_a_2;
input 	q_a_10;
input 	q_a_18;
input 	q_a_26;
input 	q_a_7;
input 	q_a_23;
input 	q_a_15;
input 	q_a_31;
input 	q_a_29;
input 	q_a_13;
input 	q_a_28;
input 	q_a_12;
input 	q_a_27;
input 	q_a_11;
input 	q_a_25;
input 	q_a_9;
input 	q_a_24;
input 	q_a_8;
input 	q_a_6;
input 	q_a_14;
input 	q_a_22;
input 	q_a_30;
input 	q_a_5;
input 	q_a_21;
input 	q_a_4;
input 	q_a_20;
input 	q_a_3;
input 	q_a_19;
input 	q_a_1;
input 	q_a_17;
input 	q_a_0;
input 	q_a_16;
input 	readdata_2;
input 	readdata_10;
input 	readdata_18;
input 	readdata_26;
input 	readdata_7;
input 	readdata_23;
input 	readdata_15;
input 	readdata_31;
input 	readdata_29;
input 	readdata_13;
input 	readdata_28;
input 	readdata_12;
input 	readdata_27;
input 	readdata_11;
input 	readdata_25;
input 	readdata_9;
input 	readdata_24;
input 	readdata_8;
input 	readdata_6;
input 	readdata_14;
input 	readdata_22;
input 	readdata_30;
input 	readdata_5;
input 	readdata_21;
input 	readdata_4;
input 	readdata_20;
input 	readdata_3;
input 	readdata_19;
input 	readdata_1;
input 	readdata_17;
input 	readdata_0;
input 	readdata_16;
input 	r_sync_rst;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
output 	hold_waitrequest;
input 	d_address_offset_field_0;
input 	d_write;
input 	d_address_tag_field_2;
input 	d_address_tag_field_1;
input 	d_address_tag_field_0;
input 	d_address_line_field_5;
input 	d_address_line_field_4;
input 	d_address_line_field_3;
input 	d_address_line_field_2;
input 	d_address_line_field_1;
input 	d_address_line_field_0;
input 	d_address_offset_field_2;
input 	d_address_offset_field_1;
output 	m0_write;
input 	d_writedata_11;
input 	d_byteenable_0;
input 	d_writedata_10;
input 	d_writedata_9;
input 	d_writedata_8;
input 	d_writedata_13;
input 	d_writedata_12;
input 	d_writedata_21;
input 	d_writedata_20;
input 	d_writedata_25;
input 	d_writedata_17;
input 	d_writedata_24;
input 	d_writedata_16;
input 	d_writedata_27;
input 	d_writedata_19;
input 	d_writedata_26;
input 	d_writedata_18;
input 	d_writedata_23;
input 	d_writedata_15;
input 	d_writedata_22;
input 	d_writedata_14;
input 	d_read;
output 	suppress_change_dest_id;
output 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
output 	saved_grant_01;
output 	mem_used_11;
output 	WideOr0;
output 	av_waitrequest;
input 	d_byteenable_1;
input 	d_writedata_2;
input 	d_writedata_0;
input 	d_writedata_3;
input 	d_writedata_1;
input 	hbreak_enabled;
input 	i_read;
output 	src0_valid;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	ic_fill_line_6;
output 	Equal1;
output 	src0_valid1;
output 	src1_valid;
output 	saved_grant_1;
output 	rf_source_valid;
output 	src1_valid1;
output 	src2_valid;
output 	saved_grant_11;
input 	d_writedata_6;
input 	d_writedata_4;
input 	d_writedata_7;
input 	d_writedata_5;
output 	WideOr1;
output 	suppress_change_dest_id1;
output 	WideOr01;
output 	WideOr02;
output 	nonposted_cmd_accepted;
input 	ic_fill_line_5;
output 	src_data_46;
output 	src_payload;
input 	ic_fill_ap_offset_0;
output 	src_data_38;
input 	ic_fill_line_1;
output 	src_data_42;
input 	ic_fill_line_0;
output 	src_data_41;
input 	ic_fill_ap_offset_2;
output 	src_data_40;
input 	ic_fill_ap_offset_1;
output 	src_data_39;
input 	ic_fill_line_4;
output 	src_data_45;
input 	ic_fill_line_3;
output 	src_data_44;
input 	ic_fill_line_2;
output 	src_data_43;
output 	src_payload1;
output 	src_data_32;
output 	src_payload2;
output 	src_payload3;
output 	WideOr11;
output 	src_data_2;
output 	src_data_10;
output 	src_data_18;
output 	src_data_26;
output 	src_data_7;
output 	src_data_23;
output 	src_data_15;
output 	src_data_31;
output 	src_data_29;
output 	src_data_13;
output 	src_data_28;
output 	src_data_12;
output 	src_data_27;
output 	src_data_11;
output 	src_data_25;
output 	src_data_9;
output 	src_data_24;
output 	src_data_8;
output 	src_data_6;
output 	src_data_14;
output 	src_data_22;
output 	src_data_30;
output 	src_data_5;
output 	src_data_21;
output 	src_data_4;
output 	src_data_20;
output 	src_data_3;
output 	src_data_19;
output 	src_data_1;
output 	src_data_17;
output 	src_data_0;
output 	src_data_16;
output 	src_payload4;
output 	src_data_51;
output 	src_data_33;
output 	src_data_110;
output 	src_data_47;
output 	src_data_210;
output 	src_data_281;
output 	src_data_311;
output 	src_data_271;
output 	src_data_291;
output 	src_data_301;
output 	src_data_01;
output 	src_data_231;
output 	src_data_261;
output 	src_data_221;
output 	src_data_241;
output 	src_data_251;
output 	src_data_161;
output 	src_data_151;
output 	src_data_131;
output 	src_data_141;
output 	src_data_121;
output 	src_data_111;
output 	src_data_81;
output 	src_payload5;
output 	src_data_381;
output 	src_data_391;
output 	src_data_401;
output 	src_data_411;
output 	src_data_421;
output 	src_data_431;
output 	src_data_441;
output 	src_data_451;
output 	src_data_461;
output 	src_data_471;
output 	src_data_321;
output 	src_payload6;
output 	src_data_331;
output 	src_payload7;
input 	d_byteenable_2;
output 	src_data_34;
output 	src_payload8;
input 	d_byteenable_3;
output 	src_data_35;
output 	src_data_191;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
input 	d_writedata_31;
output 	src_payload12;
input 	d_writedata_29;
output 	src_payload13;
output 	src_payload14;
output 	src_data_181;
input 	d_writedata_28;
output 	src_payload15;
output 	src_payload16;
output 	src_data_171;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
input 	d_writedata_30;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_data_101;
output 	src_payload29;
output 	src_payload30;
output 	src_data_91;
output 	src_payload31;
output 	src_payload32;
output 	src_payload33;
output 	src_payload34;
output 	src_payload35;
output 	src_payload36;
output 	src_data_211;
output 	src_data_201;
output 	src_data_71;
output 	src_data_61;
output 	src_payload37;
output 	src_data_351;
output 	src_payload38;
output 	src_payload39;
output 	src_data_341;
output 	src_payload40;
output 	src_payload41;
output 	src_payload42;
output 	src_payload43;
output 	src_payload44;
output 	src_payload45;
output 	src_payload46;
output 	src_payload47;
output 	src_payload48;
output 	src_payload49;
output 	src_payload50;
output 	src_payload51;
output 	src_payload52;
output 	src_payload53;
output 	src_data_332;
output 	src_payload54;
output 	src_payload55;
output 	src_payload56;
output 	src_payload57;
output 	src_payload58;
output 	src_payload59;
output 	src_payload60;
output 	src_payload61;
output 	src_payload62;
output 	src_payload63;
output 	src_payload64;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ad9833_comp_0_avalon_slave_0_agent_rsp_fifo|mem_used[1]~q ;
wire \router|always1~0_combout ;
wire \router|always1~1_combout ;
wire \ad9833_comp_0_avalon_slave_0_agent|m0_write~1_combout ;
wire \ad9833_comp_0_avalon_slave_0_translator|av_waitrequest_generated~0_combout ;
wire \ad9833_comp_0_avalon_slave_0_translator|read_latency_shift_reg[0]~q ;
wire \router|Equal2~0_combout ;
wire \cmd_demux|src2_valid~0_combout ;
wire \nios2_qsys_0_data_master_limiter|has_pending_responses~q ;
wire \nios2_qsys_0_data_master_limiter|last_dest_id[0]~q ;
wire \nios2_qsys_0_data_master_limiter|last_channel[2]~q ;
wire \ad9833_comp_0_avalon_slave_0_translator|read_latency_shift_reg~0_combout ;
wire \nios2_qsys_0_data_master_agent|cp_valid~0_combout ;
wire \nios2_qsys_0_jtag_debug_module_translator|read_latency_shift_reg[0]~q ;
wire \nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][71]~q ;
wire \nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][53]~q ;
wire \rsp_demux_001|src0_valid~0_combout ;
wire \onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][71]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][53]~q ;
wire \rsp_demux_002|src0_valid~0_combout ;
wire \ad9833_comp_0_avalon_slave_0_agent_rsp_fifo|mem[0][58]~q ;
wire \nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][58]~q ;
wire \onchip_memory2_0_s1_agent_rsp_fifo|mem[0][58]~q ;
wire \nios2_qsys_0_instruction_master_limiter|last_dest_id[0]~q ;
wire \nios2_qsys_0_instruction_master_limiter|has_pending_responses~q ;
wire \nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|write~0_combout ;
wire \nios2_qsys_0_instruction_master_limiter|last_dest_id[1]~q ;
wire \onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ;
wire \onchip_memory2_0_s1_agent|rf_source_valid~0_combout ;
wire \onchip_memory2_0_s1_translator|read_latency_shift_reg~1_combout ;
wire \rsp_demux_001|src1_valid~0_combout ;
wire \rsp_demux_002|src1_valid~0_combout ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[2]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[10]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[18]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[26]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[7]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[23]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[15]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[31]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[29]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[13]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[28]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[12]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[27]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[11]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[25]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[9]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[24]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[8]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[6]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[14]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[22]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[30]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[5]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[21]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[4]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[20]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[3]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[19]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[1]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[17]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[0]~q ;
wire \nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[16]~q ;


embedded_system_embedded_system_mm_interconnect_0_router_001 router_001(
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.ic_fill_line_6(ic_fill_line_6),
	.Equal1(Equal1));

embedded_system_embedded_system_mm_interconnect_0_router router(
	.d_address_tag_field_2(d_address_tag_field_2),
	.d_address_tag_field_1(d_address_tag_field_1),
	.d_address_tag_field_0(d_address_tag_field_0),
	.d_address_line_field_5(d_address_line_field_5),
	.d_address_line_field_4(d_address_line_field_4),
	.d_address_line_field_3(d_address_line_field_3),
	.always1(\router|always1~0_combout ),
	.d_address_line_field_2(d_address_line_field_2),
	.d_address_line_field_1(d_address_line_field_1),
	.d_address_line_field_0(d_address_line_field_0),
	.d_address_offset_field_2(d_address_offset_field_2),
	.d_address_offset_field_1(d_address_offset_field_1),
	.always11(\router|always1~1_combout ),
	.Equal2(\router|Equal2~0_combout ));

embedded_system_altera_avalon_sc_fifo_2 onchip_memory2_0_s1_agent_rsp_fifo(
	.reset(r_sync_rst),
	.hold_waitrequest(hold_waitrequest),
	.d_read(d_read),
	.saved_grant_0(saved_grant_01),
	.mem_used_1(mem_used_11),
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_71_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][71]~q ),
	.mem_53_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][53]~q ),
	.mem_58_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][58]~q ),
	.i_read(i_read),
	.saved_grant_1(saved_grant_11),
	.rf_source_valid(\onchip_memory2_0_s1_agent|rf_source_valid~0_combout ),
	.read_latency_shift_reg(\onchip_memory2_0_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

embedded_system_altera_merlin_slave_agent_2 onchip_memory2_0_s1_agent(
	.d_read(d_read),
	.saved_grant_0(saved_grant_01),
	.i_read(i_read),
	.src1_valid(src1_valid1),
	.src2_valid(src2_valid),
	.saved_grant_1(saved_grant_11),
	.rf_source_valid(\onchip_memory2_0_s1_agent|rf_source_valid~0_combout ));

embedded_system_altera_avalon_sc_fifo_1 nios2_qsys_0_jtag_debug_module_agent_rsp_fifo(
	.reset(r_sync_rst),
	.d_read(d_read),
	.saved_grant_0(saved_grant_0),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_1),
	.read_latency_shift_reg_0(\nios2_qsys_0_jtag_debug_module_translator|read_latency_shift_reg[0]~q ),
	.mem_71_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][71]~q ),
	.mem_53_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][53]~q ),
	.mem_58_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][58]~q ),
	.i_read(i_read),
	.write(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(saved_grant_1),
	.rf_source_valid(rf_source_valid),
	.clk(clk_clk));

embedded_system_altera_merlin_slave_agent_1 nios2_qsys_0_jtag_debug_module_agent(
	.d_read(d_read),
	.saved_grant_0(saved_grant_0),
	.i_read(i_read),
	.src0_valid(src0_valid1),
	.src1_valid(src1_valid),
	.saved_grant_1(saved_grant_1),
	.rf_source_valid(rf_source_valid));

embedded_system_altera_avalon_sc_fifo ad9833_comp_0_avalon_slave_0_agent_rsp_fifo(
	.reset(r_sync_rst),
	.mem_used_1(\ad9833_comp_0_avalon_slave_0_agent_rsp_fifo|mem_used[1]~q ),
	.m0_write(\ad9833_comp_0_avalon_slave_0_agent|m0_write~1_combout ),
	.av_waitrequest_generated(\ad9833_comp_0_avalon_slave_0_translator|av_waitrequest_generated~0_combout ),
	.d_read(d_read),
	.read_latency_shift_reg_0(\ad9833_comp_0_avalon_slave_0_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg(\ad9833_comp_0_avalon_slave_0_translator|read_latency_shift_reg~0_combout ),
	.mem_58_0(\ad9833_comp_0_avalon_slave_0_agent_rsp_fifo|mem[0][58]~q ),
	.clk(clk_clk));

embedded_system_altera_merlin_slave_agent ad9833_comp_0_avalon_slave_0_agent(
	.mem_used_1(\ad9833_comp_0_avalon_slave_0_agent_rsp_fifo|mem_used[1]~q ),
	.hold_waitrequest(hold_waitrequest),
	.d_address_offset_field_0(d_address_offset_field_0),
	.d_write(d_write),
	.always1(\router|always1~0_combout ),
	.always11(\router|always1~1_combout ),
	.m0_write(m0_write),
	.m0_write1(\ad9833_comp_0_avalon_slave_0_agent|m0_write~1_combout ));

embedded_system_altera_merlin_master_agent nios2_qsys_0_data_master_agent(
	.r_sync_rst(r_sync_rst),
	.hold_waitrequest1(hold_waitrequest),
	.d_write(d_write),
	.d_read(d_read),
	.suppress_change_dest_id(suppress_change_dest_id),
	.WideOr0(WideOr0),
	.av_waitrequest1(av_waitrequest),
	.cp_valid(\nios2_qsys_0_data_master_agent|cp_valid~0_combout ),
	.clk(clk_clk));

embedded_system_altera_merlin_slave_translator_2 onchip_memory2_0_s1_translator(
	.reset(r_sync_rst),
	.hold_waitrequest(hold_waitrequest),
	.mem_used_1(mem_used_11),
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg(\onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ),
	.rf_source_valid(\onchip_memory2_0_s1_agent|rf_source_valid~0_combout ),
	.read_latency_shift_reg1(\onchip_memory2_0_s1_translator|read_latency_shift_reg~1_combout ),
	.clk(clk_clk));

embedded_system_altera_merlin_slave_translator_1 nios2_qsys_0_jtag_debug_module_translator(
	.av_readdata({readdata_31,readdata_30,readdata_29,readdata_28,readdata_27,readdata_26,readdata_25,readdata_24,readdata_23,readdata_22,readdata_21,readdata_20,readdata_19,readdata_18,readdata_17,readdata_16,readdata_15,readdata_14,readdata_13,readdata_12,readdata_11,readdata_10,readdata_9,
readdata_8,readdata_7,readdata_6,readdata_5,readdata_4,readdata_3,readdata_2,readdata_1,readdata_0}),
	.reset(r_sync_rst),
	.hold_waitrequest(hold_waitrequest),
	.read_latency_shift_reg_0(\nios2_qsys_0_jtag_debug_module_translator|read_latency_shift_reg[0]~q ),
	.write(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|write~0_combout ),
	.rf_source_valid(rf_source_valid),
	.av_readdata_pre_2(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_10(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_18(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_26(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_7(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_23(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_15(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_31(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_29(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_13(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_28(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_12(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_27(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_11(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_25(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_9(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_24(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_8(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_6(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_14(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_22(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_30(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_5(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_21(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_4(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_20(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_3(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_19(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_1(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_17(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_0(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_16(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[16]~q ),
	.clk(clk_clk));

embedded_system_altera_merlin_slave_translator ad9833_comp_0_avalon_slave_0_translator(
	.reset(r_sync_rst),
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.m0_write(m0_write),
	.av_waitrequest_generated(\ad9833_comp_0_avalon_slave_0_translator|av_waitrequest_generated~0_combout ),
	.d_read(d_read),
	.read_latency_shift_reg_0(\ad9833_comp_0_avalon_slave_0_translator|read_latency_shift_reg[0]~q ),
	.read_latency_shift_reg(\ad9833_comp_0_avalon_slave_0_translator|read_latency_shift_reg~0_combout ),
	.clk(clk_clk));

embedded_system_embedded_system_mm_interconnect_0_rsp_mux_001 rsp_mux_001(
	.q_a_2(q_a_2),
	.q_a_10(q_a_10),
	.q_a_18(q_a_18),
	.q_a_26(q_a_26),
	.q_a_7(q_a_7),
	.q_a_23(q_a_23),
	.q_a_15(q_a_15),
	.q_a_31(q_a_31),
	.q_a_29(q_a_29),
	.q_a_13(q_a_13),
	.q_a_28(q_a_28),
	.q_a_12(q_a_12),
	.q_a_27(q_a_27),
	.q_a_11(q_a_11),
	.q_a_25(q_a_25),
	.q_a_9(q_a_9),
	.q_a_24(q_a_24),
	.q_a_8(q_a_8),
	.q_a_6(q_a_6),
	.q_a_14(q_a_14),
	.q_a_22(q_a_22),
	.q_a_30(q_a_30),
	.q_a_5(q_a_5),
	.q_a_21(q_a_21),
	.q_a_4(q_a_4),
	.q_a_20(q_a_20),
	.q_a_3(q_a_3),
	.q_a_19(q_a_19),
	.q_a_1(q_a_1),
	.q_a_17(q_a_17),
	.q_a_0(q_a_0),
	.q_a_16(q_a_16),
	.src1_valid(\rsp_demux_001|src1_valid~0_combout ),
	.src1_valid1(\rsp_demux_002|src1_valid~0_combout ),
	.WideOr11(WideOr11),
	.av_readdata_pre_2(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[2]~q ),
	.av_readdata_pre_10(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[10]~q ),
	.av_readdata_pre_18(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[18]~q ),
	.av_readdata_pre_26(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[26]~q ),
	.av_readdata_pre_7(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[7]~q ),
	.av_readdata_pre_23(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[23]~q ),
	.av_readdata_pre_15(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[15]~q ),
	.av_readdata_pre_31(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[31]~q ),
	.av_readdata_pre_29(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[29]~q ),
	.av_readdata_pre_13(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[13]~q ),
	.av_readdata_pre_28(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[28]~q ),
	.av_readdata_pre_12(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[12]~q ),
	.av_readdata_pre_27(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[27]~q ),
	.av_readdata_pre_11(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[11]~q ),
	.av_readdata_pre_25(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[25]~q ),
	.av_readdata_pre_9(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[9]~q ),
	.av_readdata_pre_24(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[24]~q ),
	.av_readdata_pre_8(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[8]~q ),
	.av_readdata_pre_6(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[6]~q ),
	.av_readdata_pre_14(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[14]~q ),
	.av_readdata_pre_22(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[22]~q ),
	.av_readdata_pre_30(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[30]~q ),
	.av_readdata_pre_5(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[5]~q ),
	.av_readdata_pre_21(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[21]~q ),
	.av_readdata_pre_4(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[4]~q ),
	.av_readdata_pre_20(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[20]~q ),
	.av_readdata_pre_3(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[3]~q ),
	.av_readdata_pre_19(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[19]~q ),
	.av_readdata_pre_1(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[1]~q ),
	.av_readdata_pre_17(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[17]~q ),
	.av_readdata_pre_0(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[0]~q ),
	.av_readdata_pre_16(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[16]~q ),
	.src_data_5(src_data_51),
	.src_data_3(src_data_33),
	.src_data_1(src_data_110),
	.src_data_4(src_data_47),
	.src_data_2(src_data_210),
	.src_data_28(src_data_281),
	.src_data_31(src_data_311),
	.src_data_27(src_data_271),
	.src_data_29(src_data_291),
	.src_data_30(src_data_301),
	.src_data_0(src_data_01),
	.src_data_23(src_data_231),
	.src_data_26(src_data_261),
	.src_data_22(src_data_221),
	.src_data_24(src_data_241),
	.src_data_25(src_data_251),
	.src_data_16(src_data_161),
	.src_data_15(src_data_151),
	.src_data_13(src_data_131),
	.src_data_14(src_data_141),
	.src_data_12(src_data_121),
	.src_data_11(src_data_111),
	.src_data_8(src_data_81),
	.src_data_19(src_data_191),
	.src_data_18(src_data_181),
	.src_data_17(src_data_171),
	.src_data_10(src_data_101),
	.src_data_9(src_data_91),
	.src_data_21(src_data_211),
	.src_data_20(src_data_201),
	.src_data_7(src_data_71),
	.src_data_6(src_data_61));

embedded_system_embedded_system_mm_interconnect_0_rsp_mux rsp_mux(
	.q_a_2(q_a_2),
	.q_a_10(q_a_10),
	.q_a_18(q_a_18),
	.q_a_26(q_a_26),
	.q_a_7(q_a_7),
	.q_a_23(q_a_23),
	.q_a_15(q_a_15),
	.q_a_31(q_a_31),
	.q_a_29(q_a_29),
	.q_a_13(q_a_13),
	.q_a_28(q_a_28),
	.q_a_12(q_a_12),
	.q_a_27(q_a_27),
	.q_a_11(q_a_11),
	.q_a_25(q_a_25),
	.q_a_9(q_a_9),
	.q_a_24(q_a_24),
	.q_a_8(q_a_8),
	.q_a_6(q_a_6),
	.q_a_14(q_a_14),
	.q_a_22(q_a_22),
	.q_a_30(q_a_30),
	.q_a_5(q_a_5),
	.q_a_21(q_a_21),
	.q_a_4(q_a_4),
	.q_a_20(q_a_20),
	.q_a_3(q_a_3),
	.q_a_19(q_a_19),
	.q_a_1(q_a_1),
	.q_a_17(q_a_17),
	.q_a_0(q_a_0),
	.q_a_16(q_a_16),
	.hold_waitrequest(hold_waitrequest),
	.read_latency_shift_reg_0(\ad9833_comp_0_avalon_slave_0_translator|read_latency_shift_reg[0]~q ),
	.src0_valid(\rsp_demux_001|src0_valid~0_combout ),
	.src0_valid1(\rsp_demux_002|src0_valid~0_combout ),
	.WideOr11(WideOr1),
	.av_readdata_pre_2(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[2]~q ),
	.src_data_2(src_data_2),
	.av_readdata_pre_10(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[10]~q ),
	.src_data_10(src_data_10),
	.av_readdata_pre_18(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[18]~q ),
	.src_data_18(src_data_18),
	.av_readdata_pre_26(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[26]~q ),
	.src_data_26(src_data_26),
	.av_readdata_pre_7(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[7]~q ),
	.src_data_7(src_data_7),
	.av_readdata_pre_23(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[23]~q ),
	.src_data_23(src_data_23),
	.av_readdata_pre_15(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[15]~q ),
	.src_data_15(src_data_15),
	.av_readdata_pre_31(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[31]~q ),
	.src_data_31(src_data_31),
	.av_readdata_pre_29(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[29]~q ),
	.src_data_29(src_data_29),
	.av_readdata_pre_13(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[13]~q ),
	.src_data_13(src_data_13),
	.av_readdata_pre_28(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[28]~q ),
	.src_data_28(src_data_28),
	.av_readdata_pre_12(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[12]~q ),
	.src_data_12(src_data_12),
	.av_readdata_pre_27(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[27]~q ),
	.src_data_27(src_data_27),
	.av_readdata_pre_11(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[11]~q ),
	.src_data_11(src_data_11),
	.av_readdata_pre_25(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[25]~q ),
	.src_data_25(src_data_25),
	.av_readdata_pre_9(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[9]~q ),
	.src_data_9(src_data_9),
	.av_readdata_pre_24(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[24]~q ),
	.src_data_24(src_data_24),
	.av_readdata_pre_8(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[8]~q ),
	.src_data_8(src_data_8),
	.av_readdata_pre_6(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[6]~q ),
	.src_data_6(src_data_6),
	.av_readdata_pre_14(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[14]~q ),
	.src_data_14(src_data_14),
	.av_readdata_pre_22(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[22]~q ),
	.src_data_22(src_data_22),
	.av_readdata_pre_30(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[30]~q ),
	.src_data_30(src_data_30),
	.av_readdata_pre_5(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[5]~q ),
	.src_data_5(src_data_5),
	.av_readdata_pre_21(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[21]~q ),
	.src_data_21(src_data_21),
	.av_readdata_pre_4(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[4]~q ),
	.src_data_4(src_data_4),
	.av_readdata_pre_20(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[20]~q ),
	.src_data_20(src_data_20),
	.av_readdata_pre_3(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[3]~q ),
	.src_data_3(src_data_3),
	.av_readdata_pre_19(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[19]~q ),
	.src_data_19(src_data_19),
	.av_readdata_pre_1(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[1]~q ),
	.src_data_1(src_data_1),
	.av_readdata_pre_17(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[17]~q ),
	.src_data_17(src_data_17),
	.av_readdata_pre_0(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[0]~q ),
	.src_data_0(src_data_0),
	.av_readdata_pre_16(\nios2_qsys_0_jtag_debug_module_translator|av_readdata_pre[16]~q ),
	.src_data_16(src_data_16));

embedded_system_embedded_system_mm_interconnect_0_rsp_demux_001_1 rsp_demux_002(
	.read_latency_shift_reg_0(\onchip_memory2_0_s1_translator|read_latency_shift_reg[0]~q ),
	.mem_71_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][71]~q ),
	.mem_53_0(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][53]~q ),
	.src0_valid(\rsp_demux_002|src0_valid~0_combout ),
	.src1_valid(\rsp_demux_002|src1_valid~0_combout ));

embedded_system_embedded_system_mm_interconnect_0_rsp_demux_001 rsp_demux_001(
	.read_latency_shift_reg_0(\nios2_qsys_0_jtag_debug_module_translator|read_latency_shift_reg[0]~q ),
	.mem_71_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][71]~q ),
	.mem_53_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][53]~q ),
	.src0_valid(\rsp_demux_001|src0_valid~0_combout ),
	.src1_valid(\rsp_demux_001|src1_valid~0_combout ));

embedded_system_embedded_system_mm_interconnect_0_cmd_mux_001_1 cmd_mux_002(
	.r_sync_rst(r_sync_rst),
	.d_address_offset_field_0(d_address_offset_field_0),
	.d_address_tag_field_0(d_address_tag_field_0),
	.d_address_line_field_5(d_address_line_field_5),
	.d_address_line_field_4(d_address_line_field_4),
	.d_address_line_field_3(d_address_line_field_3),
	.d_address_line_field_2(d_address_line_field_2),
	.d_address_line_field_1(d_address_line_field_1),
	.d_address_line_field_0(d_address_line_field_0),
	.d_address_offset_field_2(d_address_offset_field_2),
	.d_address_offset_field_1(d_address_offset_field_1),
	.d_writedata_11(d_writedata_11),
	.d_byteenable_0(d_byteenable_0),
	.d_writedata_10(d_writedata_10),
	.d_writedata_9(d_writedata_9),
	.d_writedata_8(d_writedata_8),
	.d_writedata_13(d_writedata_13),
	.d_writedata_12(d_writedata_12),
	.d_writedata_21(d_writedata_21),
	.d_writedata_20(d_writedata_20),
	.d_writedata_25(d_writedata_25),
	.d_writedata_17(d_writedata_17),
	.d_writedata_24(d_writedata_24),
	.d_writedata_16(d_writedata_16),
	.d_writedata_27(d_writedata_27),
	.d_writedata_19(d_writedata_19),
	.d_writedata_26(d_writedata_26),
	.d_writedata_18(d_writedata_18),
	.d_writedata_23(d_writedata_23),
	.d_writedata_15(d_writedata_15),
	.d_writedata_22(d_writedata_22),
	.d_writedata_14(d_writedata_14),
	.saved_grant_0(saved_grant_01),
	.d_byteenable_1(d_byteenable_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_0(d_writedata_0),
	.d_writedata_3(d_writedata_3),
	.d_writedata_1(d_writedata_1),
	.ic_fill_line_6(ic_fill_line_6),
	.src1_valid(src1_valid1),
	.src2_valid(src2_valid),
	.read_latency_shift_reg(\onchip_memory2_0_s1_translator|read_latency_shift_reg~0_combout ),
	.saved_grant_1(saved_grant_11),
	.d_writedata_6(d_writedata_6),
	.d_writedata_4(d_writedata_4),
	.d_writedata_7(d_writedata_7),
	.d_writedata_5(d_writedata_5),
	.ic_fill_line_5(ic_fill_line_5),
	.ic_fill_ap_offset_0(ic_fill_ap_offset_0),
	.ic_fill_line_1(ic_fill_line_1),
	.ic_fill_line_0(ic_fill_line_0),
	.ic_fill_ap_offset_2(ic_fill_ap_offset_2),
	.ic_fill_ap_offset_1(ic_fill_ap_offset_1),
	.ic_fill_line_4(ic_fill_line_4),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_2(ic_fill_line_2),
	.src_payload(src_payload5),
	.src_data_38(src_data_381),
	.src_data_39(src_data_391),
	.src_data_40(src_data_401),
	.src_data_41(src_data_411),
	.src_data_42(src_data_421),
	.src_data_43(src_data_431),
	.src_data_44(src_data_441),
	.src_data_45(src_data_451),
	.src_data_46(src_data_461),
	.src_data_47(src_data_471),
	.src_data_32(src_data_321),
	.src_payload1(src_payload6),
	.src_data_33(src_data_331),
	.src_payload2(src_payload7),
	.d_byteenable_2(d_byteenable_2),
	.src_data_34(src_data_34),
	.src_payload3(src_payload8),
	.d_byteenable_3(d_byteenable_3),
	.src_data_35(src_data_35),
	.src_payload4(src_payload9),
	.src_payload5(src_payload10),
	.src_payload6(src_payload11),
	.d_writedata_31(d_writedata_31),
	.src_payload7(src_payload12),
	.d_writedata_29(d_writedata_29),
	.src_payload8(src_payload13),
	.src_payload9(src_payload14),
	.d_writedata_28(d_writedata_28),
	.src_payload10(src_payload15),
	.src_payload11(src_payload16),
	.src_payload12(src_payload17),
	.src_payload13(src_payload18),
	.src_payload14(src_payload19),
	.src_payload15(src_payload20),
	.src_payload16(src_payload21),
	.src_payload17(src_payload22),
	.src_payload18(src_payload23),
	.src_payload19(src_payload24),
	.src_payload20(src_payload25),
	.d_writedata_30(d_writedata_30),
	.src_payload21(src_payload26),
	.src_payload22(src_payload27),
	.src_payload23(src_payload28),
	.src_payload24(src_payload29),
	.src_payload25(src_payload30),
	.src_payload26(src_payload31),
	.src_payload27(src_payload32),
	.src_payload28(src_payload33),
	.src_payload29(src_payload34),
	.src_payload30(src_payload35),
	.src_payload31(src_payload36),
	.clk_clk(clk_clk));

embedded_system_embedded_system_mm_interconnect_0_cmd_mux_001 cmd_mux_001(
	.r_sync_rst(r_sync_rst),
	.d_address_offset_field_0(d_address_offset_field_0),
	.d_address_line_field_5(d_address_line_field_5),
	.d_address_line_field_4(d_address_line_field_4),
	.d_address_line_field_3(d_address_line_field_3),
	.d_address_line_field_2(d_address_line_field_2),
	.d_address_line_field_1(d_address_line_field_1),
	.d_address_line_field_0(d_address_line_field_0),
	.d_address_offset_field_2(d_address_offset_field_2),
	.d_address_offset_field_1(d_address_offset_field_1),
	.d_writedata_11(d_writedata_11),
	.d_byteenable_0(d_byteenable_0),
	.d_writedata_10(d_writedata_10),
	.d_writedata_9(d_writedata_9),
	.d_writedata_8(d_writedata_8),
	.d_writedata_13(d_writedata_13),
	.d_writedata_12(d_writedata_12),
	.d_writedata_21(d_writedata_21),
	.d_writedata_20(d_writedata_20),
	.d_writedata_25(d_writedata_25),
	.d_writedata_17(d_writedata_17),
	.d_writedata_24(d_writedata_24),
	.d_writedata_16(d_writedata_16),
	.d_writedata_27(d_writedata_27),
	.d_writedata_19(d_writedata_19),
	.d_writedata_26(d_writedata_26),
	.d_writedata_18(d_writedata_18),
	.d_writedata_23(d_writedata_23),
	.d_writedata_15(d_writedata_15),
	.d_writedata_22(d_writedata_22),
	.d_writedata_14(d_writedata_14),
	.saved_grant_0(saved_grant_0),
	.d_byteenable_1(d_byteenable_1),
	.d_writedata_2(d_writedata_2),
	.d_writedata_0(d_writedata_0),
	.d_writedata_3(d_writedata_3),
	.d_writedata_1(d_writedata_1),
	.hbreak_enabled(hbreak_enabled),
	.src0_valid(src0_valid1),
	.src1_valid(src1_valid),
	.write(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|write~0_combout ),
	.saved_grant_1(saved_grant_1),
	.d_writedata_6(d_writedata_6),
	.d_writedata_4(d_writedata_4),
	.d_writedata_7(d_writedata_7),
	.d_writedata_5(d_writedata_5),
	.ic_fill_line_5(ic_fill_line_5),
	.src_data_46(src_data_46),
	.src_payload(src_payload),
	.ic_fill_ap_offset_0(ic_fill_ap_offset_0),
	.src_data_38(src_data_38),
	.ic_fill_line_1(ic_fill_line_1),
	.src_data_42(src_data_42),
	.ic_fill_line_0(ic_fill_line_0),
	.src_data_41(src_data_41),
	.ic_fill_ap_offset_2(ic_fill_ap_offset_2),
	.src_data_40(src_data_40),
	.ic_fill_ap_offset_1(ic_fill_ap_offset_1),
	.src_data_39(src_data_39),
	.ic_fill_line_4(ic_fill_line_4),
	.src_data_45(src_data_45),
	.ic_fill_line_3(ic_fill_line_3),
	.src_data_44(src_data_44),
	.ic_fill_line_2(ic_fill_line_2),
	.src_data_43(src_data_43),
	.src_payload1(src_payload1),
	.src_data_32(src_data_32),
	.src_payload2(src_payload2),
	.src_payload3(src_payload3),
	.src_payload4(src_payload4),
	.d_byteenable_2(d_byteenable_2),
	.d_byteenable_3(d_byteenable_3),
	.d_writedata_31(d_writedata_31),
	.d_writedata_29(d_writedata_29),
	.d_writedata_28(d_writedata_28),
	.d_writedata_30(d_writedata_30),
	.src_payload5(src_payload37),
	.src_data_35(src_data_351),
	.src_payload6(src_payload38),
	.src_payload7(src_payload39),
	.src_data_34(src_data_341),
	.src_payload8(src_payload40),
	.src_payload9(src_payload41),
	.src_payload10(src_payload42),
	.src_payload11(src_payload43),
	.src_payload12(src_payload44),
	.src_payload13(src_payload45),
	.src_payload14(src_payload46),
	.src_payload15(src_payload47),
	.src_payload16(src_payload48),
	.src_payload17(src_payload49),
	.src_payload18(src_payload50),
	.src_payload19(src_payload51),
	.src_payload20(src_payload52),
	.src_payload21(src_payload53),
	.src_data_33(src_data_332),
	.src_payload22(src_payload54),
	.src_payload23(src_payload55),
	.src_payload24(src_payload56),
	.src_payload25(src_payload57),
	.src_payload26(src_payload58),
	.src_payload27(src_payload59),
	.src_payload28(src_payload60),
	.src_payload29(src_payload61),
	.src_payload30(src_payload62),
	.src_payload31(src_payload63),
	.src_payload32(src_payload64),
	.clk_clk(clk_clk));

embedded_system_embedded_system_mm_interconnect_0_cmd_demux_001 cmd_demux_001(
	.hold_waitrequest(hold_waitrequest),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_1),
	.mem_used_11(mem_used_11),
	.last_dest_id_0(\nios2_qsys_0_instruction_master_limiter|last_dest_id[0]~q ),
	.has_pending_responses(\nios2_qsys_0_instruction_master_limiter|has_pending_responses~q ),
	.i_read(i_read),
	.src0_valid(src0_valid),
	.Equal1(Equal1),
	.src0_valid1(src0_valid1),
	.saved_grant_1(saved_grant_1),
	.last_dest_id_1(\nios2_qsys_0_instruction_master_limiter|last_dest_id[1]~q ),
	.src1_valid(src1_valid1),
	.saved_grant_11(saved_grant_11),
	.WideOr0(WideOr01),
	.WideOr01(WideOr02));

embedded_system_embedded_system_mm_interconnect_0_cmd_demux cmd_demux(
	.wait_latency_counter_1(wait_latency_counter_1),
	.wait_latency_counter_0(wait_latency_counter_0),
	.hold_waitrequest(hold_waitrequest),
	.d_address_offset_field_0(d_address_offset_field_0),
	.d_write(d_write),
	.d_address_tag_field_2(d_address_tag_field_2),
	.d_address_tag_field_1(d_address_tag_field_1),
	.d_address_tag_field_0(d_address_tag_field_0),
	.always1(\router|always1~0_combout ),
	.always11(\router|always1~1_combout ),
	.m0_write(m0_write),
	.d_read(d_read),
	.Equal2(\router|Equal2~0_combout ),
	.src2_valid(\cmd_demux|src2_valid~0_combout ),
	.has_pending_responses(\nios2_qsys_0_data_master_limiter|has_pending_responses~q ),
	.last_dest_id_0(\nios2_qsys_0_data_master_limiter|last_dest_id[0]~q ),
	.last_channel_2(\nios2_qsys_0_data_master_limiter|last_channel[2]~q ),
	.saved_grant_0(saved_grant_0),
	.waitrequest(waitrequest),
	.mem_used_1(mem_used_1),
	.saved_grant_01(saved_grant_01),
	.mem_used_11(mem_used_11),
	.WideOr01(WideOr0),
	.cp_valid(\nios2_qsys_0_data_master_agent|cp_valid~0_combout ),
	.src1_valid(src1_valid),
	.src2_valid1(src2_valid));

embedded_system_altera_merlin_traffic_limiter_1 nios2_qsys_0_instruction_master_limiter(
	.reset(r_sync_rst),
	.mem_58_0(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][58]~q ),
	.mem_58_01(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][58]~q ),
	.last_dest_id_0(\nios2_qsys_0_instruction_master_limiter|last_dest_id[0]~q ),
	.has_pending_responses1(\nios2_qsys_0_instruction_master_limiter|has_pending_responses~q ),
	.src0_valid(src0_valid),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.ic_fill_line_6(ic_fill_line_6),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,Equal1,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd}),
	.last_dest_id_1(\nios2_qsys_0_instruction_master_limiter|last_dest_id[1]~q ),
	.suppress_change_dest_id(suppress_change_dest_id1),
	.WideOr0(WideOr01),
	.WideOr01(WideOr02),
	.nonposted_cmd_accepted1(nonposted_cmd_accepted),
	.src1_valid(\rsp_demux_001|src1_valid~0_combout ),
	.src1_valid1(\rsp_demux_002|src1_valid~0_combout ),
	.clk(clk_clk));

embedded_system_altera_merlin_traffic_limiter nios2_qsys_0_data_master_limiter(
	.reset(r_sync_rst),
	.d_write(d_write),
	.d_address_tag_field_2(d_address_tag_field_2),
	.d_address_tag_field_1(d_address_tag_field_1),
	.d_address_tag_field_0(d_address_tag_field_0),
	.read_latency_shift_reg_0(\ad9833_comp_0_avalon_slave_0_translator|read_latency_shift_reg[0]~q ),
	.cmd_sink_data({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\router|Equal2~0_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd}),
	.cmd_sink_channel({\cmd_demux|src2_valid~0_combout ,gnd,gnd}),
	.has_pending_responses1(\nios2_qsys_0_data_master_limiter|has_pending_responses~q ),
	.last_dest_id_0(\nios2_qsys_0_data_master_limiter|last_dest_id[0]~q ),
	.last_channel_2(\nios2_qsys_0_data_master_limiter|last_channel[2]~q ),
	.suppress_change_dest_id(suppress_change_dest_id),
	.WideOr0(WideOr0),
	.cp_valid(\nios2_qsys_0_data_master_agent|cp_valid~0_combout ),
	.src0_valid(\rsp_demux_001|src0_valid~0_combout ),
	.src0_valid1(\rsp_demux_002|src0_valid~0_combout ),
	.mem_58_0(\ad9833_comp_0_avalon_slave_0_agent_rsp_fifo|mem[0][58]~q ),
	.mem_58_01(\nios2_qsys_0_jtag_debug_module_agent_rsp_fifo|mem[0][58]~q ),
	.mem_58_02(\onchip_memory2_0_s1_agent_rsp_fifo|mem[0][58]~q ),
	.clk(clk_clk));

endmodule

module embedded_system_altera_avalon_sc_fifo (
	reset,
	mem_used_1,
	m0_write,
	av_waitrequest_generated,
	d_read,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	mem_58_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	mem_used_1;
input 	m0_write;
input 	av_waitrequest_generated;
input 	d_read;
input 	read_latency_shift_reg_0;
input 	read_latency_shift_reg;
output 	mem_58_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~1_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][89]~q ;
wire \mem~0_combout ;
wire \mem[0][58]~1_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][58] (
	.clk(clk),
	.d(\mem[0][58]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_58_0),
	.prn(vcc));
defparam \mem[0][58] .is_wysiwyg = "true";
defparam \mem[0][58] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~1 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~1 .extended_lut = "off";
defparam \mem_used[0]~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \mem_used[0]~1 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!mem_used_1),
	.datab(!m0_write),
	.datac(!av_waitrequest_generated),
	.datad(!d_read),
	.datae(!read_latency_shift_reg_0),
	.dataf(!\mem_used[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFFFF3FFF7FFF7FFF;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][89] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][89]~q ),
	.prn(vcc));
defparam \mem[1][89] .is_wysiwyg = "true";
defparam \mem[1][89] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!\mem[1][89]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem[0][58]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(!mem_58_0),
	.datad(!\mem~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem[0][58]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem[0][58]~1 .extended_lut = "off";
defparam \mem[0][58]~1 .lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam \mem[0][58]~1 .shared_arith = "off";

endmodule

module embedded_system_altera_avalon_sc_fifo_1 (
	reset,
	d_read,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_71_0,
	mem_53_0,
	mem_58_0,
	i_read,
	write,
	saved_grant_1,
	rf_source_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_read;
input 	saved_grant_0;
input 	waitrequest;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_71_0;
output 	mem_53_0;
output 	mem_58_0;
input 	i_read;
output 	write;
input 	saved_grant_1;
input 	rf_source_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][71]~q ;
wire \mem~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][53]~q ;
wire \mem~1_combout ;
wire \mem[1][89]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][71] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_71_0),
	.prn(vcc));
defparam \mem[0][71] .is_wysiwyg = "true";
defparam \mem[0][71] .power_up = "low";

dffeas \mem[0][53] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_53_0),
	.prn(vcc));
defparam \mem[0][53] .is_wysiwyg = "true";
defparam \mem[0][53] .power_up = "low";

dffeas \mem[0][58] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_58_0),
	.prn(vcc));
defparam \mem[0][58] .is_wysiwyg = "true";
defparam \mem[0][58] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(write),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!rf_source_valid),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hBF8FFFFFBF8FFFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!rf_source_valid),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hBFBFFF3FBFBFFF3F;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][71] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][71]~q ),
	.prn(vcc));
defparam \mem[1][71] .is_wysiwyg = "true";
defparam \mem[1][71] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][71]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][53] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][53]~q ),
	.prn(vcc));
defparam \mem[1][53] .is_wysiwyg = "true";
defparam \mem[1][53] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!d_read),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!i_read),
	.datae(!saved_grant_1),
	.dataf(!\mem[1][53]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h53FFFFFFFFFFFFFF;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][89] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][89]~q ),
	.prn(vcc));
defparam \mem[1][89] .is_wysiwyg = "true";
defparam \mem[1][89] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!saved_grant_0),
	.datab(!mem_used_1),
	.datac(!saved_grant_1),
	.datad(!\mem[1][89]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \mem~2 .shared_arith = "off";

endmodule

module embedded_system_altera_avalon_sc_fifo_2 (
	reset,
	hold_waitrequest,
	d_read,
	saved_grant_0,
	mem_used_1,
	read_latency_shift_reg_0,
	mem_71_0,
	mem_53_0,
	mem_58_0,
	i_read,
	saved_grant_1,
	rf_source_valid,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	hold_waitrequest;
input 	d_read;
input 	saved_grant_0;
output 	mem_used_1;
input 	read_latency_shift_reg_0;
output 	mem_71_0;
output 	mem_53_0;
output 	mem_58_0;
input 	i_read;
input 	saved_grant_1;
input 	rf_source_valid;
input 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mem_used[0]~2_combout ;
wire \mem_used[0]~q ;
wire \mem_used[1]~0_combout ;
wire \mem[1][71]~q ;
wire \mem~0_combout ;
wire \mem_used[1]~1_combout ;
wire \mem[1][53]~q ;
wire \mem~1_combout ;
wire \mem[1][89]~q ;
wire \mem~2_combout ;


dffeas \mem_used[1] (
	.clk(clk),
	.d(\mem_used[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(mem_used_1),
	.prn(vcc));
defparam \mem_used[1] .is_wysiwyg = "true";
defparam \mem_used[1] .power_up = "low";

dffeas \mem[0][71] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_71_0),
	.prn(vcc));
defparam \mem[0][71] .is_wysiwyg = "true";
defparam \mem[0][71] .power_up = "low";

dffeas \mem[0][53] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_53_0),
	.prn(vcc));
defparam \mem[0][53] .is_wysiwyg = "true";
defparam \mem[0][53] .power_up = "low";

dffeas \mem[0][58] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\mem_used[1]~1_combout ),
	.q(mem_58_0),
	.prn(vcc));
defparam \mem[0][58] .is_wysiwyg = "true";
defparam \mem[0][58] .power_up = "low";

cyclonev_lcell_comb \mem_used[0]~2 (
	.dataa(!mem_used_1),
	.datab(!read_latency_shift_reg_0),
	.datac(!\mem_used[0]~q ),
	.datad(!read_latency_shift_reg),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[0]~2 .extended_lut = "off";
defparam \mem_used[0]~2 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \mem_used[0]~2 .shared_arith = "off";

dffeas \mem_used[0] (
	.clk(clk),
	.d(\mem_used[0]~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem_used[0]~q ),
	.prn(vcc));
defparam \mem_used[0] .is_wysiwyg = "true";
defparam \mem_used[0] .power_up = "low";

cyclonev_lcell_comb \mem_used[1]~0 (
	.dataa(!hold_waitrequest),
	.datab(!mem_used_1),
	.datac(!rf_source_valid),
	.datad(!read_latency_shift_reg_0),
	.datae(!\mem_used[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~0 .extended_lut = "off";
defparam \mem_used[1]~0 .lut_mask = 64'hFF3F7F7FFF3F7F7F;
defparam \mem_used[1]~0 .shared_arith = "off";

dffeas \mem[1][71] (
	.clk(clk),
	.d(\mem~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][71]~q ),
	.prn(vcc));
defparam \mem[1][71] .is_wysiwyg = "true";
defparam \mem[1][71] .power_up = "low";

cyclonev_lcell_comb \mem~0 (
	.dataa(!mem_used_1),
	.datab(!saved_grant_1),
	.datac(!\mem[1][71]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~0 .extended_lut = "off";
defparam \mem~0 .lut_mask = 64'h2727272727272727;
defparam \mem~0 .shared_arith = "off";

cyclonev_lcell_comb \mem_used[1]~1 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!\mem_used[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem_used[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem_used[1]~1 .extended_lut = "off";
defparam \mem_used[1]~1 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \mem_used[1]~1 .shared_arith = "off";

dffeas \mem[1][53] (
	.clk(clk),
	.d(\mem~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][53]~q ),
	.prn(vcc));
defparam \mem[1][53] .is_wysiwyg = "true";
defparam \mem[1][53] .power_up = "low";

cyclonev_lcell_comb \mem~1 (
	.dataa(!d_read),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!i_read),
	.datae(!saved_grant_1),
	.dataf(!\mem[1][53]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~1 .extended_lut = "off";
defparam \mem~1 .lut_mask = 64'h53FFFFFFFFFFFFFF;
defparam \mem~1 .shared_arith = "off";

dffeas \mem[1][89] (
	.clk(clk),
	.d(\mem~2_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\mem[1][89]~q ),
	.prn(vcc));
defparam \mem[1][89] .is_wysiwyg = "true";
defparam \mem[1][89] .power_up = "low";

cyclonev_lcell_comb \mem~2 (
	.dataa(!saved_grant_0),
	.datab(!mem_used_1),
	.datac(!saved_grant_1),
	.datad(!\mem[1][89]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\mem~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \mem~2 .extended_lut = "off";
defparam \mem~2 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \mem~2 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_master_agent (
	r_sync_rst,
	hold_waitrequest1,
	d_write,
	d_read,
	suppress_change_dest_id,
	WideOr0,
	av_waitrequest1,
	cp_valid,
	clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
output 	hold_waitrequest1;
input 	d_write;
input 	d_read;
input 	suppress_change_dest_id;
input 	WideOr0;
output 	av_waitrequest1;
output 	cp_valid;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas hold_waitrequest(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(hold_waitrequest1),
	.prn(vcc));
defparam hold_waitrequest.is_wysiwyg = "true";
defparam hold_waitrequest.power_up = "low";

cyclonev_lcell_comb av_waitrequest(
	.dataa(!hold_waitrequest1),
	.datab(!suppress_change_dest_id),
	.datac(!WideOr0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest1),
	.sumout(),
	.cout(),
	.shareout());
defparam av_waitrequest.extended_lut = "off";
defparam av_waitrequest.lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam av_waitrequest.shared_arith = "off";

cyclonev_lcell_comb \cp_valid~0 (
	.dataa(!hold_waitrequest1),
	.datab(!d_write),
	.datac(!d_read),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(cp_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \cp_valid~0 .extended_lut = "off";
defparam \cp_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \cp_valid~0 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_slave_agent (
	mem_used_1,
	hold_waitrequest,
	d_address_offset_field_0,
	d_write,
	always1,
	always11,
	m0_write,
	m0_write1)/* synthesis synthesis_greybox=1 */;
input 	mem_used_1;
input 	hold_waitrequest;
input 	d_address_offset_field_0;
input 	d_write;
input 	always1;
input 	always11;
output 	m0_write;
output 	m0_write1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \m0_write~0 (
	.dataa(!mem_used_1),
	.datab(!hold_waitrequest),
	.datac(!d_address_offset_field_0),
	.datad(!d_write),
	.datae(!always1),
	.dataf(!always11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~0 .extended_lut = "off";
defparam \m0_write~0 .lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam \m0_write~0 .shared_arith = "off";

cyclonev_lcell_comb \m0_write~1 (
	.dataa(!hold_waitrequest),
	.datab(!d_address_offset_field_0),
	.datac(!d_write),
	.datad(!always1),
	.datae(!always11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(m0_write1),
	.sumout(),
	.cout(),
	.shareout());
defparam \m0_write~1 .extended_lut = "off";
defparam \m0_write~1 .lut_mask = 64'hDFFFFFFFDFFFFFFF;
defparam \m0_write~1 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_slave_agent_1 (
	d_read,
	saved_grant_0,
	i_read,
	src0_valid,
	src1_valid,
	saved_grant_1,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	d_read;
input 	saved_grant_0;
input 	i_read;
input 	src0_valid;
input 	src1_valid;
input 	saved_grant_1;
output 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!d_read),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!src0_valid),
	.datae(!src1_valid),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \rf_source_valid~0 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_slave_agent_2 (
	d_read,
	saved_grant_0,
	i_read,
	src1_valid,
	src2_valid,
	saved_grant_1,
	rf_source_valid)/* synthesis synthesis_greybox=1 */;
input 	d_read;
input 	saved_grant_0;
input 	i_read;
input 	src1_valid;
input 	src2_valid;
input 	saved_grant_1;
output 	rf_source_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \rf_source_valid~0 (
	.dataa(!d_read),
	.datab(!saved_grant_0),
	.datac(!i_read),
	.datad(!src1_valid),
	.datae(!src2_valid),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(rf_source_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_source_valid~0 .extended_lut = "off";
defparam \rf_source_valid~0 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \rf_source_valid~0 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_slave_translator (
	reset,
	wait_latency_counter_1,
	wait_latency_counter_0,
	m0_write,
	av_waitrequest_generated,
	d_read,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
output 	wait_latency_counter_1;
output 	wait_latency_counter_0;
input 	m0_write;
output 	av_waitrequest_generated;
input 	d_read;
output 	read_latency_shift_reg_0;
output 	read_latency_shift_reg;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wait_latency_counter~0_combout ;
wire \wait_latency_counter~1_combout ;


dffeas \wait_latency_counter[1] (
	.clk(clk),
	.d(\wait_latency_counter~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_1),
	.prn(vcc));
defparam \wait_latency_counter[1] .is_wysiwyg = "true";
defparam \wait_latency_counter[1] .power_up = "low";

dffeas \wait_latency_counter[0] (
	.clk(clk),
	.d(\wait_latency_counter~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(wait_latency_counter_0),
	.prn(vcc));
defparam \wait_latency_counter[0] .is_wysiwyg = "true";
defparam \wait_latency_counter[0] .power_up = "low";

cyclonev_lcell_comb \av_waitrequest_generated~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(av_waitrequest_generated),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_waitrequest_generated~0 .extended_lut = "off";
defparam \av_waitrequest_generated~0 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \av_waitrequest_generated~0 .shared_arith = "off";

dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!m0_write),
	.datab(!av_waitrequest_generated),
	.datac(!d_read),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~0 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~0 .extended_lut = "off";
defparam \wait_latency_counter~0 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \wait_latency_counter~0 .shared_arith = "off";

cyclonev_lcell_comb \wait_latency_counter~1 (
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_latency_counter~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_latency_counter~1 .extended_lut = "off";
defparam \wait_latency_counter~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \wait_latency_counter~1 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_slave_translator_1 (
	av_readdata,
	reset,
	hold_waitrequest,
	read_latency_shift_reg_0,
	write,
	rf_source_valid,
	av_readdata_pre_2,
	av_readdata_pre_10,
	av_readdata_pre_18,
	av_readdata_pre_26,
	av_readdata_pre_7,
	av_readdata_pre_23,
	av_readdata_pre_15,
	av_readdata_pre_31,
	av_readdata_pre_29,
	av_readdata_pre_13,
	av_readdata_pre_28,
	av_readdata_pre_12,
	av_readdata_pre_27,
	av_readdata_pre_11,
	av_readdata_pre_25,
	av_readdata_pre_9,
	av_readdata_pre_24,
	av_readdata_pre_8,
	av_readdata_pre_6,
	av_readdata_pre_14,
	av_readdata_pre_22,
	av_readdata_pre_30,
	av_readdata_pre_5,
	av_readdata_pre_21,
	av_readdata_pre_4,
	av_readdata_pre_20,
	av_readdata_pre_3,
	av_readdata_pre_19,
	av_readdata_pre_1,
	av_readdata_pre_17,
	av_readdata_pre_0,
	av_readdata_pre_16,
	clk)/* synthesis synthesis_greybox=1 */;
input 	[31:0] av_readdata;
input 	reset;
input 	hold_waitrequest;
output 	read_latency_shift_reg_0;
input 	write;
input 	rf_source_valid;
output 	av_readdata_pre_2;
output 	av_readdata_pre_10;
output 	av_readdata_pre_18;
output 	av_readdata_pre_26;
output 	av_readdata_pre_7;
output 	av_readdata_pre_23;
output 	av_readdata_pre_15;
output 	av_readdata_pre_31;
output 	av_readdata_pre_29;
output 	av_readdata_pre_13;
output 	av_readdata_pre_28;
output 	av_readdata_pre_12;
output 	av_readdata_pre_27;
output 	av_readdata_pre_11;
output 	av_readdata_pre_25;
output 	av_readdata_pre_9;
output 	av_readdata_pre_24;
output 	av_readdata_pre_8;
output 	av_readdata_pre_6;
output 	av_readdata_pre_14;
output 	av_readdata_pre_22;
output 	av_readdata_pre_30;
output 	av_readdata_pre_5;
output 	av_readdata_pre_21;
output 	av_readdata_pre_4;
output 	av_readdata_pre_20;
output 	av_readdata_pre_3;
output 	av_readdata_pre_19;
output 	av_readdata_pre_1;
output 	av_readdata_pre_17;
output 	av_readdata_pre_0;
output 	av_readdata_pre_16;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \read_latency_shift_reg~0_combout ;


dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(\read_latency_shift_reg~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

dffeas \av_readdata_pre[2] (
	.clk(clk),
	.d(av_readdata[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_2),
	.prn(vcc));
defparam \av_readdata_pre[2] .is_wysiwyg = "true";
defparam \av_readdata_pre[2] .power_up = "low";

dffeas \av_readdata_pre[10] (
	.clk(clk),
	.d(av_readdata[10]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_10),
	.prn(vcc));
defparam \av_readdata_pre[10] .is_wysiwyg = "true";
defparam \av_readdata_pre[10] .power_up = "low";

dffeas \av_readdata_pre[18] (
	.clk(clk),
	.d(av_readdata[18]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_18),
	.prn(vcc));
defparam \av_readdata_pre[18] .is_wysiwyg = "true";
defparam \av_readdata_pre[18] .power_up = "low";

dffeas \av_readdata_pre[26] (
	.clk(clk),
	.d(av_readdata[26]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_26),
	.prn(vcc));
defparam \av_readdata_pre[26] .is_wysiwyg = "true";
defparam \av_readdata_pre[26] .power_up = "low";

dffeas \av_readdata_pre[7] (
	.clk(clk),
	.d(av_readdata[7]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_7),
	.prn(vcc));
defparam \av_readdata_pre[7] .is_wysiwyg = "true";
defparam \av_readdata_pre[7] .power_up = "low";

dffeas \av_readdata_pre[23] (
	.clk(clk),
	.d(av_readdata[23]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_23),
	.prn(vcc));
defparam \av_readdata_pre[23] .is_wysiwyg = "true";
defparam \av_readdata_pre[23] .power_up = "low";

dffeas \av_readdata_pre[15] (
	.clk(clk),
	.d(av_readdata[15]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_15),
	.prn(vcc));
defparam \av_readdata_pre[15] .is_wysiwyg = "true";
defparam \av_readdata_pre[15] .power_up = "low";

dffeas \av_readdata_pre[31] (
	.clk(clk),
	.d(av_readdata[31]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_31),
	.prn(vcc));
defparam \av_readdata_pre[31] .is_wysiwyg = "true";
defparam \av_readdata_pre[31] .power_up = "low";

dffeas \av_readdata_pre[29] (
	.clk(clk),
	.d(av_readdata[29]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_29),
	.prn(vcc));
defparam \av_readdata_pre[29] .is_wysiwyg = "true";
defparam \av_readdata_pre[29] .power_up = "low";

dffeas \av_readdata_pre[13] (
	.clk(clk),
	.d(av_readdata[13]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_13),
	.prn(vcc));
defparam \av_readdata_pre[13] .is_wysiwyg = "true";
defparam \av_readdata_pre[13] .power_up = "low";

dffeas \av_readdata_pre[28] (
	.clk(clk),
	.d(av_readdata[28]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_28),
	.prn(vcc));
defparam \av_readdata_pre[28] .is_wysiwyg = "true";
defparam \av_readdata_pre[28] .power_up = "low";

dffeas \av_readdata_pre[12] (
	.clk(clk),
	.d(av_readdata[12]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_12),
	.prn(vcc));
defparam \av_readdata_pre[12] .is_wysiwyg = "true";
defparam \av_readdata_pre[12] .power_up = "low";

dffeas \av_readdata_pre[27] (
	.clk(clk),
	.d(av_readdata[27]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_27),
	.prn(vcc));
defparam \av_readdata_pre[27] .is_wysiwyg = "true";
defparam \av_readdata_pre[27] .power_up = "low";

dffeas \av_readdata_pre[11] (
	.clk(clk),
	.d(av_readdata[11]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_11),
	.prn(vcc));
defparam \av_readdata_pre[11] .is_wysiwyg = "true";
defparam \av_readdata_pre[11] .power_up = "low";

dffeas \av_readdata_pre[25] (
	.clk(clk),
	.d(av_readdata[25]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_25),
	.prn(vcc));
defparam \av_readdata_pre[25] .is_wysiwyg = "true";
defparam \av_readdata_pre[25] .power_up = "low";

dffeas \av_readdata_pre[9] (
	.clk(clk),
	.d(av_readdata[9]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_9),
	.prn(vcc));
defparam \av_readdata_pre[9] .is_wysiwyg = "true";
defparam \av_readdata_pre[9] .power_up = "low";

dffeas \av_readdata_pre[24] (
	.clk(clk),
	.d(av_readdata[24]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_24),
	.prn(vcc));
defparam \av_readdata_pre[24] .is_wysiwyg = "true";
defparam \av_readdata_pre[24] .power_up = "low";

dffeas \av_readdata_pre[8] (
	.clk(clk),
	.d(av_readdata[8]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_8),
	.prn(vcc));
defparam \av_readdata_pre[8] .is_wysiwyg = "true";
defparam \av_readdata_pre[8] .power_up = "low";

dffeas \av_readdata_pre[6] (
	.clk(clk),
	.d(av_readdata[6]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_6),
	.prn(vcc));
defparam \av_readdata_pre[6] .is_wysiwyg = "true";
defparam \av_readdata_pre[6] .power_up = "low";

dffeas \av_readdata_pre[14] (
	.clk(clk),
	.d(av_readdata[14]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_14),
	.prn(vcc));
defparam \av_readdata_pre[14] .is_wysiwyg = "true";
defparam \av_readdata_pre[14] .power_up = "low";

dffeas \av_readdata_pre[22] (
	.clk(clk),
	.d(av_readdata[22]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_22),
	.prn(vcc));
defparam \av_readdata_pre[22] .is_wysiwyg = "true";
defparam \av_readdata_pre[22] .power_up = "low";

dffeas \av_readdata_pre[30] (
	.clk(clk),
	.d(av_readdata[30]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_30),
	.prn(vcc));
defparam \av_readdata_pre[30] .is_wysiwyg = "true";
defparam \av_readdata_pre[30] .power_up = "low";

dffeas \av_readdata_pre[5] (
	.clk(clk),
	.d(av_readdata[5]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_5),
	.prn(vcc));
defparam \av_readdata_pre[5] .is_wysiwyg = "true";
defparam \av_readdata_pre[5] .power_up = "low";

dffeas \av_readdata_pre[21] (
	.clk(clk),
	.d(av_readdata[21]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_21),
	.prn(vcc));
defparam \av_readdata_pre[21] .is_wysiwyg = "true";
defparam \av_readdata_pre[21] .power_up = "low";

dffeas \av_readdata_pre[4] (
	.clk(clk),
	.d(av_readdata[4]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_4),
	.prn(vcc));
defparam \av_readdata_pre[4] .is_wysiwyg = "true";
defparam \av_readdata_pre[4] .power_up = "low";

dffeas \av_readdata_pre[20] (
	.clk(clk),
	.d(av_readdata[20]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_20),
	.prn(vcc));
defparam \av_readdata_pre[20] .is_wysiwyg = "true";
defparam \av_readdata_pre[20] .power_up = "low";

dffeas \av_readdata_pre[3] (
	.clk(clk),
	.d(av_readdata[3]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_3),
	.prn(vcc));
defparam \av_readdata_pre[3] .is_wysiwyg = "true";
defparam \av_readdata_pre[3] .power_up = "low";

dffeas \av_readdata_pre[19] (
	.clk(clk),
	.d(av_readdata[19]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_19),
	.prn(vcc));
defparam \av_readdata_pre[19] .is_wysiwyg = "true";
defparam \av_readdata_pre[19] .power_up = "low";

dffeas \av_readdata_pre[1] (
	.clk(clk),
	.d(av_readdata[1]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_1),
	.prn(vcc));
defparam \av_readdata_pre[1] .is_wysiwyg = "true";
defparam \av_readdata_pre[1] .power_up = "low";

dffeas \av_readdata_pre[17] (
	.clk(clk),
	.d(av_readdata[17]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_17),
	.prn(vcc));
defparam \av_readdata_pre[17] .is_wysiwyg = "true";
defparam \av_readdata_pre[17] .power_up = "low";

dffeas \av_readdata_pre[0] (
	.clk(clk),
	.d(av_readdata[0]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_0),
	.prn(vcc));
defparam \av_readdata_pre[0] .is_wysiwyg = "true";
defparam \av_readdata_pre[0] .power_up = "low";

dffeas \av_readdata_pre[16] (
	.clk(clk),
	.d(av_readdata[16]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(av_readdata_pre_16),
	.prn(vcc));
defparam \av_readdata_pre[16] .is_wysiwyg = "true";
defparam \av_readdata_pre[16] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!hold_waitrequest),
	.datab(!write),
	.datac(!rf_source_valid),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read_latency_shift_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_slave_translator_2 (
	reset,
	hold_waitrequest,
	mem_used_1,
	read_latency_shift_reg_0,
	read_latency_shift_reg,
	rf_source_valid,
	read_latency_shift_reg1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	hold_waitrequest;
input 	mem_used_1;
output 	read_latency_shift_reg_0;
output 	read_latency_shift_reg;
input 	rf_source_valid;
output 	read_latency_shift_reg1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \read_latency_shift_reg[0] (
	.clk(clk),
	.d(read_latency_shift_reg1),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(read_latency_shift_reg_0),
	.prn(vcc));
defparam \read_latency_shift_reg[0] .is_wysiwyg = "true";
defparam \read_latency_shift_reg[0] .power_up = "low";

cyclonev_lcell_comb \read_latency_shift_reg~0 (
	.dataa(!hold_waitrequest),
	.datab(!mem_used_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~0 .extended_lut = "off";
defparam \read_latency_shift_reg~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \read_latency_shift_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \read_latency_shift_reg~1 (
	.dataa(!read_latency_shift_reg),
	.datab(!rf_source_valid),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(read_latency_shift_reg1),
	.sumout(),
	.cout(),
	.shareout());
defparam \read_latency_shift_reg~1 .extended_lut = "off";
defparam \read_latency_shift_reg~1 .lut_mask = 64'h7777777777777777;
defparam \read_latency_shift_reg~1 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_traffic_limiter (
	reset,
	d_write,
	d_address_tag_field_2,
	d_address_tag_field_1,
	d_address_tag_field_0,
	read_latency_shift_reg_0,
	cmd_sink_data,
	cmd_sink_channel,
	has_pending_responses1,
	last_dest_id_0,
	last_channel_2,
	suppress_change_dest_id,
	WideOr0,
	cp_valid,
	src0_valid,
	src0_valid1,
	mem_58_0,
	mem_58_01,
	mem_58_02,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	d_write;
input 	d_address_tag_field_2;
input 	d_address_tag_field_1;
input 	d_address_tag_field_0;
input 	read_latency_shift_reg_0;
input 	[87:0] cmd_sink_data;
input 	[2:0] cmd_sink_channel;
output 	has_pending_responses1;
output 	last_dest_id_0;
output 	last_channel_2;
output 	suppress_change_dest_id;
input 	WideOr0;
input 	cp_valid;
input 	src0_valid;
input 	src0_valid1;
input 	mem_58_0;
input 	mem_58_01;
input 	mem_58_02;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \save_dest_id~0_combout ;
wire \response_sink_accepted~0_combout ;
wire \pending_response_count[0]~0_combout ;
wire \pending_response_count[0]~q ;
wire \has_pending_responses~0_combout ;


dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

dffeas \last_dest_id[0] (
	.clk(clk),
	.d(cmd_sink_data[73]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_dest_id_0),
	.prn(vcc));
defparam \last_dest_id[0] .is_wysiwyg = "true";
defparam \last_dest_id[0] .power_up = "low";

dffeas \last_channel[2] (
	.clk(clk),
	.d(cmd_sink_channel[2]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_channel_2),
	.prn(vcc));
defparam \last_channel[2] .is_wysiwyg = "true";
defparam \last_channel[2] .power_up = "low";

cyclonev_lcell_comb \suppress_change_dest_id~0 (
	.dataa(!d_write),
	.datab(!cmd_sink_channel[2]),
	.datac(!has_pending_responses1),
	.datad(!\Equal0~0_combout ),
	.datae(!last_channel_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(suppress_change_dest_id),
	.sumout(),
	.cout(),
	.shareout());
defparam \suppress_change_dest_id~0 .extended_lut = "off";
defparam \suppress_change_dest_id~0 .lut_mask = 64'hBFFFEFFFBFFFEFFF;
defparam \suppress_change_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!d_address_tag_field_2),
	.datab(!d_address_tag_field_1),
	.datac(!d_address_tag_field_0),
	.datad(!last_dest_id_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h6996699669966996;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!d_write),
	.datab(!cmd_sink_channel[2]),
	.datac(!has_pending_responses1),
	.datad(!\Equal0~0_combout ),
	.datae(!last_channel_2),
	.dataf(!cp_valid),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\save_dest_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'hFFFBFFFEFFFFFFFF;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(!mem_58_0),
	.datae(!mem_58_01),
	.dataf(!mem_58_02),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~0 (
	.dataa(!WideOr0),
	.datab(!\save_dest_id~0_combout ),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~0 .extended_lut = "off";
defparam \pending_response_count[0]~0 .lut_mask = 64'h6996699669966996;
defparam \pending_response_count[0]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!has_pending_responses1),
	.datab(!WideOr0),
	.datac(!\save_dest_id~0_combout ),
	.datad(!\pending_response_count[0]~q ),
	.datae(!\response_sink_accepted~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \has_pending_responses~0 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_traffic_limiter_1 (
	reset,
	mem_58_0,
	mem_58_01,
	last_dest_id_0,
	has_pending_responses1,
	src0_valid,
	ic_fill_tag_1,
	ic_fill_tag_0,
	ic_fill_line_6,
	cmd_sink_data,
	last_dest_id_1,
	suppress_change_dest_id,
	WideOr0,
	WideOr01,
	nonposted_cmd_accepted1,
	src1_valid,
	src1_valid1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	mem_58_0;
input 	mem_58_01;
output 	last_dest_id_0;
output 	has_pending_responses1;
input 	src0_valid;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	ic_fill_line_6;
input 	[87:0] cmd_sink_data;
output 	last_dest_id_1;
output 	suppress_change_dest_id;
input 	WideOr0;
input 	WideOr01;
output 	nonposted_cmd_accepted1;
input 	src1_valid;
input 	src1_valid1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \save_dest_id~0_combout ;
wire \response_sink_accepted~0_combout ;
wire \pending_response_count[0]~0_combout ;
wire \pending_response_count[0]~q ;
wire \has_pending_responses~0_combout ;
wire \last_dest_id[1]~0_combout ;


dffeas \last_dest_id[0] (
	.clk(clk),
	.d(cmd_sink_data[73]),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_dest_id_0),
	.prn(vcc));
defparam \last_dest_id[0] .is_wysiwyg = "true";
defparam \last_dest_id[0] .power_up = "low";

dffeas has_pending_responses(
	.clk(clk),
	.d(\has_pending_responses~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(has_pending_responses1),
	.prn(vcc));
defparam has_pending_responses.is_wysiwyg = "true";
defparam has_pending_responses.power_up = "low";

dffeas \last_dest_id[1] (
	.clk(clk),
	.d(\last_dest_id[1]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\save_dest_id~0_combout ),
	.q(last_dest_id_1),
	.prn(vcc));
defparam \last_dest_id[1] .is_wysiwyg = "true";
defparam \last_dest_id[1] .power_up = "low";

cyclonev_lcell_comb \suppress_change_dest_id~0 (
	.dataa(!last_dest_id_0),
	.datab(!has_pending_responses1),
	.datac(!ic_fill_tag_1),
	.datad(!ic_fill_tag_0),
	.datae(!ic_fill_line_6),
	.dataf(!last_dest_id_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(suppress_change_dest_id),
	.sumout(),
	.cout(),
	.shareout());
defparam \suppress_change_dest_id~0 .extended_lut = "off";
defparam \suppress_change_dest_id~0 .lut_mask = 64'hB77B7BB77BB7B77B;
defparam \suppress_change_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb nonposted_cmd_accepted(
	.dataa(!src0_valid),
	.datab(!cmd_sink_data[73]),
	.datac(!suppress_change_dest_id),
	.datad(!WideOr0),
	.datae(!WideOr01),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(nonposted_cmd_accepted1),
	.sumout(),
	.cout(),
	.shareout());
defparam nonposted_cmd_accepted.extended_lut = "off";
defparam nonposted_cmd_accepted.lut_mask = 64'hD1FFFFFFD1FFFFFF;
defparam nonposted_cmd_accepted.shared_arith = "off";

cyclonev_lcell_comb \save_dest_id~0 (
	.dataa(!src0_valid),
	.datab(!suppress_change_dest_id),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\save_dest_id~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \save_dest_id~0 .extended_lut = "off";
defparam \save_dest_id~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \save_dest_id~0 .shared_arith = "off";

cyclonev_lcell_comb \response_sink_accepted~0 (
	.dataa(!mem_58_0),
	.datab(!mem_58_01),
	.datac(!src1_valid),
	.datad(!src1_valid1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\response_sink_accepted~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \response_sink_accepted~0 .extended_lut = "off";
defparam \response_sink_accepted~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \response_sink_accepted~0 .shared_arith = "off";

cyclonev_lcell_comb \pending_response_count[0]~0 (
	.dataa(!nonposted_cmd_accepted1),
	.datab(!\pending_response_count[0]~q ),
	.datac(!\response_sink_accepted~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\pending_response_count[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \pending_response_count[0]~0 .extended_lut = "off";
defparam \pending_response_count[0]~0 .lut_mask = 64'h9696969696969696;
defparam \pending_response_count[0]~0 .shared_arith = "off";

dffeas \pending_response_count[0] (
	.clk(clk),
	.d(\pending_response_count[0]~0_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\pending_response_count[0]~q ),
	.prn(vcc));
defparam \pending_response_count[0] .is_wysiwyg = "true";
defparam \pending_response_count[0] .power_up = "low";

cyclonev_lcell_comb \has_pending_responses~0 (
	.dataa(!has_pending_responses1),
	.datab(!nonposted_cmd_accepted1),
	.datac(!\pending_response_count[0]~q ),
	.datad(!\response_sink_accepted~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\has_pending_responses~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \has_pending_responses~0 .extended_lut = "off";
defparam \has_pending_responses~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \has_pending_responses~0 .shared_arith = "off";

cyclonev_lcell_comb \last_dest_id[1]~0 (
	.dataa(!cmd_sink_data[73]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\last_dest_id[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \last_dest_id[1]~0 .extended_lut = "off";
defparam \last_dest_id[1]~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \last_dest_id[1]~0 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_mm_interconnect_0_cmd_demux (
	wait_latency_counter_1,
	wait_latency_counter_0,
	hold_waitrequest,
	d_address_offset_field_0,
	d_write,
	d_address_tag_field_2,
	d_address_tag_field_1,
	d_address_tag_field_0,
	always1,
	always11,
	m0_write,
	d_read,
	Equal2,
	src2_valid,
	has_pending_responses,
	last_dest_id_0,
	last_channel_2,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	saved_grant_01,
	mem_used_11,
	WideOr01,
	cp_valid,
	src1_valid,
	src2_valid1)/* synthesis synthesis_greybox=1 */;
input 	wait_latency_counter_1;
input 	wait_latency_counter_0;
input 	hold_waitrequest;
input 	d_address_offset_field_0;
input 	d_write;
input 	d_address_tag_field_2;
input 	d_address_tag_field_1;
input 	d_address_tag_field_0;
input 	always1;
input 	always11;
input 	m0_write;
input 	d_read;
input 	Equal2;
output 	src2_valid;
input 	has_pending_responses;
input 	last_dest_id_0;
input 	last_channel_2;
input 	saved_grant_0;
input 	waitrequest;
input 	mem_used_1;
input 	saved_grant_01;
input 	mem_used_11;
output 	WideOr01;
input 	cp_valid;
output 	src1_valid;
output 	src2_valid1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sink_ready~0_combout ;
wire \sink_ready~1_combout ;
wire \src2_valid~1_combout ;


cyclonev_lcell_comb \src2_valid~0 (
	.dataa(!d_address_offset_field_0),
	.datab(!d_write),
	.datac(!always1),
	.datad(!always11),
	.datae(!Equal2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~0 .extended_lut = "off";
defparam \src2_valid~0 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \src2_valid~0 .shared_arith = "off";

cyclonev_lcell_comb WideOr0(
	.dataa(!wait_latency_counter_1),
	.datab(!wait_latency_counter_0),
	.datac(!m0_write),
	.datad(!src2_valid),
	.datae(!\sink_ready~0_combout ),
	.dataf(!\sink_ready~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr0.extended_lut = "off";
defparam WideOr0.lut_mask = 64'hFFFFFFFFFFFFFFF7;
defparam WideOr0.shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!d_write),
	.datab(!Equal2),
	.datac(!has_pending_responses),
	.datad(!last_dest_id_0),
	.datae(!cp_valid),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~2 (
	.dataa(!d_address_offset_field_0),
	.datab(!d_write),
	.datac(!always1),
	.datad(!always11),
	.datae(!Equal2),
	.dataf(!\src2_valid~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src2_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~2 .extended_lut = "off";
defparam \src2_valid~2 .lut_mask = 64'hFFFFFFFDFFFFFFFF;
defparam \src2_valid~2 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~0 (
	.dataa(!d_address_tag_field_2),
	.datab(!d_address_tag_field_1),
	.datac(!d_address_tag_field_0),
	.datad(!saved_grant_0),
	.datae(!waitrequest),
	.dataf(!mem_used_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~0 .extended_lut = "off";
defparam \sink_ready~0 .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \sink_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \sink_ready~1 (
	.dataa(!hold_waitrequest),
	.datab(!saved_grant_01),
	.datac(!mem_used_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sink_ready~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sink_ready~1 .extended_lut = "off";
defparam \sink_ready~1 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \sink_ready~1 .shared_arith = "off";

cyclonev_lcell_comb \src2_valid~1 (
	.dataa(!hold_waitrequest),
	.datab(!d_write),
	.datac(!d_read),
	.datad(!has_pending_responses),
	.datae(!last_channel_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src2_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src2_valid~1 .extended_lut = "off";
defparam \src2_valid~1 .lut_mask = 64'hFF7FFFFFFF7FFFFF;
defparam \src2_valid~1 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_mm_interconnect_0_cmd_demux_001 (
	hold_waitrequest,
	waitrequest,
	mem_used_1,
	mem_used_11,
	last_dest_id_0,
	has_pending_responses,
	i_read,
	src0_valid,
	Equal1,
	src0_valid1,
	saved_grant_1,
	last_dest_id_1,
	src1_valid,
	saved_grant_11,
	WideOr0,
	WideOr01)/* synthesis synthesis_greybox=1 */;
input 	hold_waitrequest;
input 	waitrequest;
input 	mem_used_1;
input 	mem_used_11;
input 	last_dest_id_0;
input 	has_pending_responses;
input 	i_read;
output 	src0_valid;
input 	Equal1;
output 	src0_valid1;
input 	saved_grant_1;
input 	last_dest_id_1;
output 	src1_valid;
input 	saved_grant_11;
output 	WideOr0;
output 	WideOr01;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!hold_waitrequest),
	.datab(!i_read),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'h7777777777777777;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src0_valid~1 (
	.dataa(!last_dest_id_0),
	.datab(!has_pending_responses),
	.datac(!src0_valid),
	.datad(!Equal1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~1 .extended_lut = "off";
defparam \src0_valid~1 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \src0_valid~1 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!has_pending_responses),
	.datab(!src0_valid),
	.datac(!Equal1),
	.datad(!last_dest_id_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \src1_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr0),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~0 .extended_lut = "off";
defparam \WideOr0~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \WideOr0~0 .shared_arith = "off";

cyclonev_lcell_comb \WideOr0~1 (
	.dataa(!hold_waitrequest),
	.datab(!mem_used_11),
	.datac(!saved_grant_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr01),
	.sumout(),
	.cout(),
	.shareout());
defparam \WideOr0~1 .extended_lut = "off";
defparam \WideOr0~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \WideOr0~1 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_mm_interconnect_0_cmd_mux_001 (
	r_sync_rst,
	d_address_offset_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	d_address_line_field_2,
	d_address_line_field_1,
	d_address_line_field_0,
	d_address_offset_field_2,
	d_address_offset_field_1,
	d_writedata_11,
	d_byteenable_0,
	d_writedata_10,
	d_writedata_9,
	d_writedata_8,
	d_writedata_13,
	d_writedata_12,
	d_writedata_21,
	d_writedata_20,
	d_writedata_25,
	d_writedata_17,
	d_writedata_24,
	d_writedata_16,
	d_writedata_27,
	d_writedata_19,
	d_writedata_26,
	d_writedata_18,
	d_writedata_23,
	d_writedata_15,
	d_writedata_22,
	d_writedata_14,
	saved_grant_0,
	d_byteenable_1,
	d_writedata_2,
	d_writedata_0,
	d_writedata_3,
	d_writedata_1,
	hbreak_enabled,
	src0_valid,
	src1_valid,
	write,
	saved_grant_1,
	d_writedata_6,
	d_writedata_4,
	d_writedata_7,
	d_writedata_5,
	ic_fill_line_5,
	src_data_46,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	ic_fill_line_1,
	src_data_42,
	ic_fill_line_0,
	src_data_41,
	ic_fill_ap_offset_2,
	src_data_40,
	ic_fill_ap_offset_1,
	src_data_39,
	ic_fill_line_4,
	src_data_45,
	ic_fill_line_3,
	src_data_44,
	ic_fill_line_2,
	src_data_43,
	src_payload1,
	src_data_32,
	src_payload2,
	src_payload3,
	src_payload4,
	d_byteenable_2,
	d_byteenable_3,
	d_writedata_31,
	d_writedata_29,
	d_writedata_28,
	d_writedata_30,
	src_payload5,
	src_data_35,
	src_payload6,
	src_payload7,
	src_data_34,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_data_33,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	d_address_offset_field_0;
input 	d_address_line_field_5;
input 	d_address_line_field_4;
input 	d_address_line_field_3;
input 	d_address_line_field_2;
input 	d_address_line_field_1;
input 	d_address_line_field_0;
input 	d_address_offset_field_2;
input 	d_address_offset_field_1;
input 	d_writedata_11;
input 	d_byteenable_0;
input 	d_writedata_10;
input 	d_writedata_9;
input 	d_writedata_8;
input 	d_writedata_13;
input 	d_writedata_12;
input 	d_writedata_21;
input 	d_writedata_20;
input 	d_writedata_25;
input 	d_writedata_17;
input 	d_writedata_24;
input 	d_writedata_16;
input 	d_writedata_27;
input 	d_writedata_19;
input 	d_writedata_26;
input 	d_writedata_18;
input 	d_writedata_23;
input 	d_writedata_15;
input 	d_writedata_22;
input 	d_writedata_14;
output 	saved_grant_0;
input 	d_byteenable_1;
input 	d_writedata_2;
input 	d_writedata_0;
input 	d_writedata_3;
input 	d_writedata_1;
input 	hbreak_enabled;
input 	src0_valid;
input 	src1_valid;
input 	write;
output 	saved_grant_1;
input 	d_writedata_6;
input 	d_writedata_4;
input 	d_writedata_7;
input 	d_writedata_5;
input 	ic_fill_line_5;
output 	src_data_46;
output 	src_payload;
input 	ic_fill_ap_offset_0;
output 	src_data_38;
input 	ic_fill_line_1;
output 	src_data_42;
input 	ic_fill_line_0;
output 	src_data_41;
input 	ic_fill_ap_offset_2;
output 	src_data_40;
input 	ic_fill_ap_offset_1;
output 	src_data_39;
input 	ic_fill_line_4;
output 	src_data_45;
input 	ic_fill_line_3;
output 	src_data_44;
input 	ic_fill_line_2;
output 	src_data_43;
output 	src_payload1;
output 	src_data_32;
output 	src_payload2;
output 	src_payload3;
output 	src_payload4;
input 	d_byteenable_2;
input 	d_byteenable_3;
input 	d_writedata_31;
input 	d_writedata_29;
input 	d_writedata_28;
input 	d_writedata_30;
output 	src_payload5;
output 	src_data_35;
output 	src_payload6;
output 	src_payload7;
output 	src_data_34;
output 	src_payload8;
output 	src_payload9;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
output 	src_payload21;
output 	src_data_33;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
output 	src_payload32;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


embedded_system_altera_merlin_arbitrator arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.src0_valid(src0_valid),
	.src1_valid(src1_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.write(write),
	.packet_in_progress(\packet_in_progress~q ),
	.saved_grant_1(saved_grant_1),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!d_address_line_field_5),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!d_address_offset_field_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!d_address_line_field_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!d_address_line_field_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!d_address_offset_field_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!d_address_offset_field_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!d_address_line_field_4),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!d_address_line_field_3),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!d_address_line_field_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!saved_grant_0),
	.datab(!hbreak_enabled),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!d_byteenable_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!d_writedata_24),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!d_writedata_20),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!d_writedata_19),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!d_writedata_16),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!d_writedata_25),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!d_writedata_26),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!d_writedata_27),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!d_writedata_21),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!d_writedata_18),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!d_writedata_17),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!d_writedata_10),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!d_byteenable_1),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!d_writedata_23),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!d_writedata_15),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!d_writedata_13),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!d_writedata_12),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!d_writedata_11),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!d_writedata_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!d_writedata_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!d_writedata_14),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~32 (
	.dataa(!d_writedata_22),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~32 .extended_lut = "off";
defparam \src_payload~32 .lut_mask = 64'h7777777777777777;
defparam \src_payload~32 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!src0_valid),
	.datad(!src1_valid),
	.datae(!\packet_in_progress~q ),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_arbitrator (
	reset,
	saved_grant_0,
	src0_valid,
	src1_valid,
	grant_0,
	write,
	packet_in_progress,
	saved_grant_1,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	src0_valid;
input 	src1_valid;
output 	grant_0;
input 	write;
input 	packet_in_progress;
input 	saved_grant_1;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!\top_priority_reg[0]~q ),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!src0_valid),
	.datad(!src1_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!\top_priority_reg[0]~q ),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!src0_valid),
	.datad(!src1_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!write),
	.datac(!src0_valid),
	.datad(!src1_valid),
	.datae(!packet_in_progress),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module embedded_system_embedded_system_mm_interconnect_0_cmd_mux_001_1 (
	r_sync_rst,
	d_address_offset_field_0,
	d_address_tag_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	d_address_line_field_2,
	d_address_line_field_1,
	d_address_line_field_0,
	d_address_offset_field_2,
	d_address_offset_field_1,
	d_writedata_11,
	d_byteenable_0,
	d_writedata_10,
	d_writedata_9,
	d_writedata_8,
	d_writedata_13,
	d_writedata_12,
	d_writedata_21,
	d_writedata_20,
	d_writedata_25,
	d_writedata_17,
	d_writedata_24,
	d_writedata_16,
	d_writedata_27,
	d_writedata_19,
	d_writedata_26,
	d_writedata_18,
	d_writedata_23,
	d_writedata_15,
	d_writedata_22,
	d_writedata_14,
	saved_grant_0,
	d_byteenable_1,
	d_writedata_2,
	d_writedata_0,
	d_writedata_3,
	d_writedata_1,
	ic_fill_line_6,
	src1_valid,
	src2_valid,
	read_latency_shift_reg,
	saved_grant_1,
	d_writedata_6,
	d_writedata_4,
	d_writedata_7,
	d_writedata_5,
	ic_fill_line_5,
	ic_fill_ap_offset_0,
	ic_fill_line_1,
	ic_fill_line_0,
	ic_fill_ap_offset_2,
	ic_fill_ap_offset_1,
	ic_fill_line_4,
	ic_fill_line_3,
	ic_fill_line_2,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_32,
	src_payload1,
	src_data_33,
	src_payload2,
	d_byteenable_2,
	src_data_34,
	src_payload3,
	d_byteenable_3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	d_writedata_31,
	src_payload7,
	d_writedata_29,
	src_payload8,
	src_payload9,
	d_writedata_28,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	d_writedata_30,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	r_sync_rst;
input 	d_address_offset_field_0;
input 	d_address_tag_field_0;
input 	d_address_line_field_5;
input 	d_address_line_field_4;
input 	d_address_line_field_3;
input 	d_address_line_field_2;
input 	d_address_line_field_1;
input 	d_address_line_field_0;
input 	d_address_offset_field_2;
input 	d_address_offset_field_1;
input 	d_writedata_11;
input 	d_byteenable_0;
input 	d_writedata_10;
input 	d_writedata_9;
input 	d_writedata_8;
input 	d_writedata_13;
input 	d_writedata_12;
input 	d_writedata_21;
input 	d_writedata_20;
input 	d_writedata_25;
input 	d_writedata_17;
input 	d_writedata_24;
input 	d_writedata_16;
input 	d_writedata_27;
input 	d_writedata_19;
input 	d_writedata_26;
input 	d_writedata_18;
input 	d_writedata_23;
input 	d_writedata_15;
input 	d_writedata_22;
input 	d_writedata_14;
output 	saved_grant_0;
input 	d_byteenable_1;
input 	d_writedata_2;
input 	d_writedata_0;
input 	d_writedata_3;
input 	d_writedata_1;
input 	ic_fill_line_6;
input 	src1_valid;
input 	src2_valid;
input 	read_latency_shift_reg;
output 	saved_grant_1;
input 	d_writedata_6;
input 	d_writedata_4;
input 	d_writedata_7;
input 	d_writedata_5;
input 	ic_fill_line_5;
input 	ic_fill_ap_offset_0;
input 	ic_fill_line_1;
input 	ic_fill_line_0;
input 	ic_fill_ap_offset_2;
input 	ic_fill_ap_offset_1;
input 	ic_fill_line_4;
input 	ic_fill_line_3;
input 	ic_fill_line_2;
output 	src_payload;
output 	src_data_38;
output 	src_data_39;
output 	src_data_40;
output 	src_data_41;
output 	src_data_42;
output 	src_data_43;
output 	src_data_44;
output 	src_data_45;
output 	src_data_46;
output 	src_data_47;
output 	src_data_32;
output 	src_payload1;
output 	src_data_33;
output 	src_payload2;
input 	d_byteenable_2;
output 	src_data_34;
output 	src_payload3;
input 	d_byteenable_3;
output 	src_data_35;
output 	src_payload4;
output 	src_payload5;
output 	src_payload6;
input 	d_writedata_31;
output 	src_payload7;
input 	d_writedata_29;
output 	src_payload8;
output 	src_payload9;
input 	d_writedata_28;
output 	src_payload10;
output 	src_payload11;
output 	src_payload12;
output 	src_payload13;
output 	src_payload14;
output 	src_payload15;
output 	src_payload16;
output 	src_payload17;
output 	src_payload18;
output 	src_payload19;
output 	src_payload20;
input 	d_writedata_30;
output 	src_payload21;
output 	src_payload22;
output 	src_payload23;
output 	src_payload24;
output 	src_payload25;
output 	src_payload26;
output 	src_payload27;
output 	src_payload28;
output 	src_payload29;
output 	src_payload30;
output 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \arb|grant[0]~0_combout ;
wire \arb|grant[1]~1_combout ;
wire \packet_in_progress~0_combout ;
wire \packet_in_progress~q ;
wire \update_grant~0_combout ;


embedded_system_altera_merlin_arbitrator_1 arb(
	.reset(r_sync_rst),
	.saved_grant_0(saved_grant_0),
	.src1_valid(src1_valid),
	.src2_valid(src2_valid),
	.grant_0(\arb|grant[0]~0_combout ),
	.read_latency_shift_reg(read_latency_shift_reg),
	.packet_in_progress(\packet_in_progress~q ),
	.saved_grant_1(saved_grant_1),
	.grant_1(\arb|grant[1]~1_combout ),
	.clk(clk_clk));

dffeas \saved_grant[0] (
	.clk(clk_clk),
	.d(\arb|grant[0]~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_0),
	.prn(vcc));
defparam \saved_grant[0] .is_wysiwyg = "true";
defparam \saved_grant[0] .power_up = "low";

dffeas \saved_grant[1] (
	.clk(clk_clk),
	.d(\arb|grant[1]~1_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_grant~0_combout ),
	.q(saved_grant_1),
	.prn(vcc));
defparam \saved_grant[1] .is_wysiwyg = "true";
defparam \saved_grant[1] .power_up = "low";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

cyclonev_lcell_comb \src_data[38] (
	.dataa(!d_address_offset_field_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_38),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[38] .extended_lut = "off";
defparam \src_data[38] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[38] .shared_arith = "off";

cyclonev_lcell_comb \src_data[39] (
	.dataa(!d_address_offset_field_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_39),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[39] .extended_lut = "off";
defparam \src_data[39] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[39] .shared_arith = "off";

cyclonev_lcell_comb \src_data[40] (
	.dataa(!d_address_offset_field_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_ap_offset_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_40),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[40] .extended_lut = "off";
defparam \src_data[40] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[40] .shared_arith = "off";

cyclonev_lcell_comb \src_data[41] (
	.dataa(!d_address_line_field_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_41),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[41] .extended_lut = "off";
defparam \src_data[41] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[41] .shared_arith = "off";

cyclonev_lcell_comb \src_data[42] (
	.dataa(!d_address_line_field_1),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_42),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[42] .extended_lut = "off";
defparam \src_data[42] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[42] .shared_arith = "off";

cyclonev_lcell_comb \src_data[43] (
	.dataa(!d_address_line_field_2),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_43),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[43] .extended_lut = "off";
defparam \src_data[43] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[43] .shared_arith = "off";

cyclonev_lcell_comb \src_data[44] (
	.dataa(!d_address_line_field_3),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_44),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[44] .extended_lut = "off";
defparam \src_data[44] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[44] .shared_arith = "off";

cyclonev_lcell_comb \src_data[45] (
	.dataa(!d_address_line_field_4),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_45),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[45] .extended_lut = "off";
defparam \src_data[45] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[45] .shared_arith = "off";

cyclonev_lcell_comb \src_data[46] (
	.dataa(!d_address_line_field_5),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(!ic_fill_line_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_46),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[46] .extended_lut = "off";
defparam \src_data[46] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[46] .shared_arith = "off";

cyclonev_lcell_comb \src_data[47] (
	.dataa(!d_address_tag_field_0),
	.datab(!saved_grant_0),
	.datac(!ic_fill_line_6),
	.datad(!saved_grant_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_47),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[47] .extended_lut = "off";
defparam \src_data[47] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[47] .shared_arith = "off";

cyclonev_lcell_comb \src_data[32] (
	.dataa(!d_byteenable_0),
	.datab(!saved_grant_0),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_32),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[32] .extended_lut = "off";
defparam \src_data[32] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[32] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~1 (
	.dataa(!d_writedata_10),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~1 .extended_lut = "off";
defparam \src_payload~1 .lut_mask = 64'h7777777777777777;
defparam \src_payload~1 .shared_arith = "off";

cyclonev_lcell_comb \src_data[33] (
	.dataa(!saved_grant_0),
	.datab(!d_byteenable_1),
	.datac(!saved_grant_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_33),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[33] .extended_lut = "off";
defparam \src_data[33] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[33] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~2 (
	.dataa(!d_writedata_18),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~2 .extended_lut = "off";
defparam \src_payload~2 .lut_mask = 64'h7777777777777777;
defparam \src_payload~2 .shared_arith = "off";

cyclonev_lcell_comb \src_data[34] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_34),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[34] .extended_lut = "off";
defparam \src_data[34] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[34] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~3 (
	.dataa(!d_writedata_26),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~3 .extended_lut = "off";
defparam \src_payload~3 .lut_mask = 64'h7777777777777777;
defparam \src_payload~3 .shared_arith = "off";

cyclonev_lcell_comb \src_data[35] (
	.dataa(!saved_grant_0),
	.datab(!saved_grant_1),
	.datac(!d_byteenable_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_35),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[35] .extended_lut = "off";
defparam \src_data[35] .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src_data[35] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~4 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~4 .extended_lut = "off";
defparam \src_payload~4 .lut_mask = 64'h7777777777777777;
defparam \src_payload~4 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~5 (
	.dataa(!d_writedata_23),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~5 .extended_lut = "off";
defparam \src_payload~5 .lut_mask = 64'h7777777777777777;
defparam \src_payload~5 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~6 (
	.dataa(!d_writedata_15),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~6 .extended_lut = "off";
defparam \src_payload~6 .lut_mask = 64'h7777777777777777;
defparam \src_payload~6 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~7 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_31),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~7 .extended_lut = "off";
defparam \src_payload~7 .lut_mask = 64'h7777777777777777;
defparam \src_payload~7 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~8 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_29),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~8 .extended_lut = "off";
defparam \src_payload~8 .lut_mask = 64'h7777777777777777;
defparam \src_payload~8 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~9 (
	.dataa(!d_writedata_13),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~9 .extended_lut = "off";
defparam \src_payload~9 .lut_mask = 64'h7777777777777777;
defparam \src_payload~9 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~10 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_28),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~10 .extended_lut = "off";
defparam \src_payload~10 .lut_mask = 64'h7777777777777777;
defparam \src_payload~10 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~11 (
	.dataa(!d_writedata_12),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~11 .extended_lut = "off";
defparam \src_payload~11 .lut_mask = 64'h7777777777777777;
defparam \src_payload~11 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~12 (
	.dataa(!d_writedata_27),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~12 .extended_lut = "off";
defparam \src_payload~12 .lut_mask = 64'h7777777777777777;
defparam \src_payload~12 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~13 (
	.dataa(!d_writedata_11),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~13 .extended_lut = "off";
defparam \src_payload~13 .lut_mask = 64'h7777777777777777;
defparam \src_payload~13 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~14 (
	.dataa(!d_writedata_25),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~14 .extended_lut = "off";
defparam \src_payload~14 .lut_mask = 64'h7777777777777777;
defparam \src_payload~14 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~15 (
	.dataa(!d_writedata_9),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~15 .extended_lut = "off";
defparam \src_payload~15 .lut_mask = 64'h7777777777777777;
defparam \src_payload~15 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~16 (
	.dataa(!d_writedata_24),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~16 .extended_lut = "off";
defparam \src_payload~16 .lut_mask = 64'h7777777777777777;
defparam \src_payload~16 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~17 (
	.dataa(!d_writedata_8),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~17 .extended_lut = "off";
defparam \src_payload~17 .lut_mask = 64'h7777777777777777;
defparam \src_payload~17 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~18 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~18 .extended_lut = "off";
defparam \src_payload~18 .lut_mask = 64'h7777777777777777;
defparam \src_payload~18 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~19 (
	.dataa(!d_writedata_14),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~19 .extended_lut = "off";
defparam \src_payload~19 .lut_mask = 64'h7777777777777777;
defparam \src_payload~19 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~20 (
	.dataa(!d_writedata_22),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~20 .extended_lut = "off";
defparam \src_payload~20 .lut_mask = 64'h7777777777777777;
defparam \src_payload~20 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~21 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_30),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~21 .extended_lut = "off";
defparam \src_payload~21 .lut_mask = 64'h7777777777777777;
defparam \src_payload~21 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~22 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~22 .extended_lut = "off";
defparam \src_payload~22 .lut_mask = 64'h7777777777777777;
defparam \src_payload~22 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~23 (
	.dataa(!d_writedata_21),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~23 .extended_lut = "off";
defparam \src_payload~23 .lut_mask = 64'h7777777777777777;
defparam \src_payload~23 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~24 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~24 .extended_lut = "off";
defparam \src_payload~24 .lut_mask = 64'h7777777777777777;
defparam \src_payload~24 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~25 (
	.dataa(!d_writedata_20),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~25 .extended_lut = "off";
defparam \src_payload~25 .lut_mask = 64'h7777777777777777;
defparam \src_payload~25 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~26 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~26 .extended_lut = "off";
defparam \src_payload~26 .lut_mask = 64'h7777777777777777;
defparam \src_payload~26 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~27 (
	.dataa(!d_writedata_19),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~27 .extended_lut = "off";
defparam \src_payload~27 .lut_mask = 64'h7777777777777777;
defparam \src_payload~27 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~28 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~28 .extended_lut = "off";
defparam \src_payload~28 .lut_mask = 64'h7777777777777777;
defparam \src_payload~28 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~29 (
	.dataa(!d_writedata_17),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~29 .extended_lut = "off";
defparam \src_payload~29 .lut_mask = 64'h7777777777777777;
defparam \src_payload~29 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~30 (
	.dataa(!saved_grant_0),
	.datab(!d_writedata_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~30 .extended_lut = "off";
defparam \src_payload~30 .lut_mask = 64'h7777777777777777;
defparam \src_payload~30 .shared_arith = "off";

cyclonev_lcell_comb \src_payload~31 (
	.dataa(!d_writedata_16),
	.datab(!saved_grant_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_payload31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~31 .extended_lut = "off";
defparam \src_payload~31 .lut_mask = 64'h7777777777777777;
defparam \src_payload~31 .shared_arith = "off";

cyclonev_lcell_comb \packet_in_progress~0 (
	.dataa(!\update_grant~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\packet_in_progress~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \packet_in_progress~0 .extended_lut = "off";
defparam \packet_in_progress~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \packet_in_progress~0 .shared_arith = "off";

dffeas packet_in_progress(
	.clk(clk_clk),
	.d(\packet_in_progress~0_combout ),
	.asdata(vcc),
	.clrn(!r_sync_rst),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\packet_in_progress~q ),
	.prn(vcc));
defparam packet_in_progress.is_wysiwyg = "true";
defparam packet_in_progress.power_up = "low";

cyclonev_lcell_comb \update_grant~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src1_valid),
	.datad(!src2_valid),
	.datae(!\packet_in_progress~q ),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_grant~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_grant~0 .extended_lut = "off";
defparam \update_grant~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \update_grant~0 .shared_arith = "off";

endmodule

module embedded_system_altera_merlin_arbitrator_1 (
	reset,
	saved_grant_0,
	src1_valid,
	src2_valid,
	grant_0,
	read_latency_shift_reg,
	packet_in_progress,
	saved_grant_1,
	grant_1,
	clk)/* synthesis synthesis_greybox=1 */;
input 	reset;
input 	saved_grant_0;
input 	src1_valid;
input 	src2_valid;
output 	grant_0;
input 	read_latency_shift_reg;
input 	packet_in_progress;
input 	saved_grant_1;
output 	grant_1;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \top_priority_reg[0]~1_combout ;
wire \top_priority_reg[0]~0_combout ;
wire \top_priority_reg[0]~q ;
wire \top_priority_reg[1]~q ;


cyclonev_lcell_comb \grant[0]~0 (
	.dataa(!\top_priority_reg[0]~q ),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!src1_valid),
	.datad(!src2_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[0]~0 .extended_lut = "off";
defparam \grant[0]~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \grant[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \grant[1]~1 (
	.dataa(!\top_priority_reg[0]~q ),
	.datab(!\top_priority_reg[1]~q ),
	.datac(!src1_valid),
	.datad(!src2_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(grant_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \grant[1]~1 .extended_lut = "off";
defparam \grant[1]~1 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \grant[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~1 (
	.dataa(!grant_1),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~1 .extended_lut = "off";
defparam \top_priority_reg[0]~1 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \top_priority_reg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \top_priority_reg[0]~0 (
	.dataa(!saved_grant_0),
	.datab(!read_latency_shift_reg),
	.datac(!src1_valid),
	.datad(!src2_valid),
	.datae(!packet_in_progress),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\top_priority_reg[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \top_priority_reg[0]~0 .extended_lut = "off";
defparam \top_priority_reg[0]~0 .lut_mask = 64'hFFFF7BB7FFFFB77B;
defparam \top_priority_reg[0]~0 .shared_arith = "off";

dffeas \top_priority_reg[0] (
	.clk(clk),
	.d(\top_priority_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[0]~q ),
	.prn(vcc));
defparam \top_priority_reg[0] .is_wysiwyg = "true";
defparam \top_priority_reg[0] .power_up = "low";

dffeas \top_priority_reg[1] (
	.clk(clk),
	.d(grant_0),
	.asdata(vcc),
	.clrn(!reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\top_priority_reg[0]~0_combout ),
	.q(\top_priority_reg[1]~q ),
	.prn(vcc));
defparam \top_priority_reg[1] .is_wysiwyg = "true";
defparam \top_priority_reg[1] .power_up = "low";

endmodule

module embedded_system_embedded_system_mm_interconnect_0_router (
	d_address_tag_field_2,
	d_address_tag_field_1,
	d_address_tag_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	always1,
	d_address_line_field_2,
	d_address_line_field_1,
	d_address_line_field_0,
	d_address_offset_field_2,
	d_address_offset_field_1,
	always11,
	Equal2)/* synthesis synthesis_greybox=1 */;
input 	d_address_tag_field_2;
input 	d_address_tag_field_1;
input 	d_address_tag_field_0;
input 	d_address_line_field_5;
input 	d_address_line_field_4;
input 	d_address_line_field_3;
output 	always1;
input 	d_address_line_field_2;
input 	d_address_line_field_1;
input 	d_address_line_field_0;
input 	d_address_offset_field_2;
input 	d_address_offset_field_1;
output 	always11;
output 	Equal2;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \always1~0 (
	.dataa(!d_address_tag_field_2),
	.datab(!d_address_tag_field_1),
	.datac(!d_address_tag_field_0),
	.datad(!d_address_line_field_5),
	.datae(!d_address_line_field_4),
	.dataf(!d_address_line_field_3),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always1),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~0 .extended_lut = "off";
defparam \always1~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \always1~0 .shared_arith = "off";

cyclonev_lcell_comb \always1~1 (
	.dataa(!d_address_line_field_2),
	.datab(!d_address_line_field_1),
	.datac(!d_address_line_field_0),
	.datad(!d_address_offset_field_2),
	.datae(!d_address_offset_field_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(always11),
	.sumout(),
	.cout(),
	.shareout());
defparam \always1~1 .extended_lut = "off";
defparam \always1~1 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \always1~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!d_address_tag_field_2),
	.datab(!d_address_tag_field_1),
	.datac(!d_address_tag_field_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal2),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \Equal2~0 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_mm_interconnect_0_router_001 (
	ic_fill_tag_1,
	ic_fill_tag_0,
	ic_fill_line_6,
	Equal1)/* synthesis synthesis_greybox=1 */;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	ic_fill_line_6;
output 	Equal1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \Equal1~0 (
	.dataa(!ic_fill_tag_1),
	.datab(!ic_fill_tag_0),
	.datac(!ic_fill_line_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal1),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal1~0 .extended_lut = "off";
defparam \Equal1~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \Equal1~0 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_mm_interconnect_0_rsp_demux_001 (
	read_latency_shift_reg_0,
	mem_71_0,
	mem_53_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_71_0;
input 	mem_53_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_71_0),
	.datac(!mem_53_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_71_0),
	.datac(!mem_53_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_mm_interconnect_0_rsp_demux_001_1 (
	read_latency_shift_reg_0,
	mem_71_0,
	mem_53_0,
	src0_valid,
	src1_valid)/* synthesis synthesis_greybox=1 */;
input 	read_latency_shift_reg_0;
input 	mem_71_0;
input 	mem_53_0;
output 	src0_valid;
output 	src1_valid;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \src0_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_71_0),
	.datac(!mem_53_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src0_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src0_valid~0 .extended_lut = "off";
defparam \src0_valid~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \src0_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \src1_valid~0 (
	.dataa(!read_latency_shift_reg_0),
	.datab(!mem_71_0),
	.datac(!mem_53_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src1_valid),
	.sumout(),
	.cout(),
	.shareout());
defparam \src1_valid~0 .extended_lut = "off";
defparam \src1_valid~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \src1_valid~0 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_mm_interconnect_0_rsp_mux (
	q_a_2,
	q_a_10,
	q_a_18,
	q_a_26,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_29,
	q_a_13,
	q_a_28,
	q_a_12,
	q_a_27,
	q_a_11,
	q_a_25,
	q_a_9,
	q_a_24,
	q_a_8,
	q_a_6,
	q_a_14,
	q_a_22,
	q_a_30,
	q_a_5,
	q_a_21,
	q_a_4,
	q_a_20,
	q_a_3,
	q_a_19,
	q_a_1,
	q_a_17,
	q_a_0,
	q_a_16,
	hold_waitrequest,
	read_latency_shift_reg_0,
	src0_valid,
	src0_valid1,
	WideOr11,
	av_readdata_pre_2,
	src_data_2,
	av_readdata_pre_10,
	src_data_10,
	av_readdata_pre_18,
	src_data_18,
	av_readdata_pre_26,
	src_data_26,
	av_readdata_pre_7,
	src_data_7,
	av_readdata_pre_23,
	src_data_23,
	av_readdata_pre_15,
	src_data_15,
	av_readdata_pre_31,
	src_data_31,
	av_readdata_pre_29,
	src_data_29,
	av_readdata_pre_13,
	src_data_13,
	av_readdata_pre_28,
	src_data_28,
	av_readdata_pre_12,
	src_data_12,
	av_readdata_pre_27,
	src_data_27,
	av_readdata_pre_11,
	src_data_11,
	av_readdata_pre_25,
	src_data_25,
	av_readdata_pre_9,
	src_data_9,
	av_readdata_pre_24,
	src_data_24,
	av_readdata_pre_8,
	src_data_8,
	av_readdata_pre_6,
	src_data_6,
	av_readdata_pre_14,
	src_data_14,
	av_readdata_pre_22,
	src_data_22,
	av_readdata_pre_30,
	src_data_30,
	av_readdata_pre_5,
	src_data_5,
	av_readdata_pre_21,
	src_data_21,
	av_readdata_pre_4,
	src_data_4,
	av_readdata_pre_20,
	src_data_20,
	av_readdata_pre_3,
	src_data_3,
	av_readdata_pre_19,
	src_data_19,
	av_readdata_pre_1,
	src_data_1,
	av_readdata_pre_17,
	src_data_17,
	av_readdata_pre_0,
	src_data_0,
	av_readdata_pre_16,
	src_data_16)/* synthesis synthesis_greybox=1 */;
input 	q_a_2;
input 	q_a_10;
input 	q_a_18;
input 	q_a_26;
input 	q_a_7;
input 	q_a_23;
input 	q_a_15;
input 	q_a_31;
input 	q_a_29;
input 	q_a_13;
input 	q_a_28;
input 	q_a_12;
input 	q_a_27;
input 	q_a_11;
input 	q_a_25;
input 	q_a_9;
input 	q_a_24;
input 	q_a_8;
input 	q_a_6;
input 	q_a_14;
input 	q_a_22;
input 	q_a_30;
input 	q_a_5;
input 	q_a_21;
input 	q_a_4;
input 	q_a_20;
input 	q_a_3;
input 	q_a_19;
input 	q_a_1;
input 	q_a_17;
input 	q_a_0;
input 	q_a_16;
input 	hold_waitrequest;
input 	read_latency_shift_reg_0;
input 	src0_valid;
input 	src0_valid1;
output 	WideOr11;
input 	av_readdata_pre_2;
output 	src_data_2;
input 	av_readdata_pre_10;
output 	src_data_10;
input 	av_readdata_pre_18;
output 	src_data_18;
input 	av_readdata_pre_26;
output 	src_data_26;
input 	av_readdata_pre_7;
output 	src_data_7;
input 	av_readdata_pre_23;
output 	src_data_23;
input 	av_readdata_pre_15;
output 	src_data_15;
input 	av_readdata_pre_31;
output 	src_data_31;
input 	av_readdata_pre_29;
output 	src_data_29;
input 	av_readdata_pre_13;
output 	src_data_13;
input 	av_readdata_pre_28;
output 	src_data_28;
input 	av_readdata_pre_12;
output 	src_data_12;
input 	av_readdata_pre_27;
output 	src_data_27;
input 	av_readdata_pre_11;
output 	src_data_11;
input 	av_readdata_pre_25;
output 	src_data_25;
input 	av_readdata_pre_9;
output 	src_data_9;
input 	av_readdata_pre_24;
output 	src_data_24;
input 	av_readdata_pre_8;
output 	src_data_8;
input 	av_readdata_pre_6;
output 	src_data_6;
input 	av_readdata_pre_14;
output 	src_data_14;
input 	av_readdata_pre_22;
output 	src_data_22;
input 	av_readdata_pre_30;
output 	src_data_30;
input 	av_readdata_pre_5;
output 	src_data_5;
input 	av_readdata_pre_21;
output 	src_data_21;
input 	av_readdata_pre_4;
output 	src_data_4;
input 	av_readdata_pre_20;
output 	src_data_20;
input 	av_readdata_pre_3;
output 	src_data_3;
input 	av_readdata_pre_19;
output 	src_data_19;
input 	av_readdata_pre_1;
output 	src_data_1;
input 	av_readdata_pre_17;
output 	src_data_17;
input 	av_readdata_pre_0;
output 	src_data_0;
input 	av_readdata_pre_16;
output 	src_data_16;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \src_payload~0_combout ;


cyclonev_lcell_comb WideOr1(
	.dataa(!read_latency_shift_reg_0),
	.datab(!src0_valid),
	.datac(!src0_valid1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[2] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_2),
	.datae(!q_a_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2] .extended_lut = "off";
defparam \src_data[2] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[2] .shared_arith = "off";

cyclonev_lcell_comb \src_data[10] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_10),
	.datae(!q_a_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10] .extended_lut = "off";
defparam \src_data[10] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[10] .shared_arith = "off";

cyclonev_lcell_comb \src_data[18] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_18),
	.datae(!q_a_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18] .extended_lut = "off";
defparam \src_data[18] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[18] .shared_arith = "off";

cyclonev_lcell_comb \src_data[26] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_26),
	.datae(!q_a_26),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26] .extended_lut = "off";
defparam \src_data[26] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[26] .shared_arith = "off";

cyclonev_lcell_comb \src_data[7] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_7),
	.datae(!q_a_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7] .extended_lut = "off";
defparam \src_data[7] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[7] .shared_arith = "off";

cyclonev_lcell_comb \src_data[23] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_23),
	.datae(!q_a_23),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23] .extended_lut = "off";
defparam \src_data[23] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[23] .shared_arith = "off";

cyclonev_lcell_comb \src_data[15] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_15),
	.datae(!q_a_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15] .extended_lut = "off";
defparam \src_data[15] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[15] .shared_arith = "off";

cyclonev_lcell_comb \src_data[31] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_31),
	.datae(!q_a_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31] .extended_lut = "off";
defparam \src_data[31] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[31] .shared_arith = "off";

cyclonev_lcell_comb \src_data[29] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_29),
	.datad(!q_a_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29] .extended_lut = "off";
defparam \src_data[29] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[29] .shared_arith = "off";

cyclonev_lcell_comb \src_data[13] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_13),
	.datad(!q_a_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13] .extended_lut = "off";
defparam \src_data[13] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[13] .shared_arith = "off";

cyclonev_lcell_comb \src_data[28] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_28),
	.datae(!q_a_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28] .extended_lut = "off";
defparam \src_data[28] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[28] .shared_arith = "off";

cyclonev_lcell_comb \src_data[12] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_12),
	.datae(!q_a_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12] .extended_lut = "off";
defparam \src_data[12] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[12] .shared_arith = "off";

cyclonev_lcell_comb \src_data[27] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_27),
	.datae(!q_a_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27] .extended_lut = "off";
defparam \src_data[27] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[27] .shared_arith = "off";

cyclonev_lcell_comb \src_data[11] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_11),
	.datae(!q_a_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11] .extended_lut = "off";
defparam \src_data[11] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[11] .shared_arith = "off";

cyclonev_lcell_comb \src_data[25] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_25),
	.datae(!q_a_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25] .extended_lut = "off";
defparam \src_data[25] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[25] .shared_arith = "off";

cyclonev_lcell_comb \src_data[9] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_9),
	.datae(!q_a_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9] .extended_lut = "off";
defparam \src_data[9] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[9] .shared_arith = "off";

cyclonev_lcell_comb \src_data[24] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_24),
	.datad(!q_a_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24] .extended_lut = "off";
defparam \src_data[24] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[24] .shared_arith = "off";

cyclonev_lcell_comb \src_data[8] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_8),
	.datad(!q_a_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8] .extended_lut = "off";
defparam \src_data[8] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[8] .shared_arith = "off";

cyclonev_lcell_comb \src_data[6] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_6),
	.datad(!q_a_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6] .extended_lut = "off";
defparam \src_data[6] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[6] .shared_arith = "off";

cyclonev_lcell_comb \src_data[14] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_14),
	.datae(!q_a_14),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14] .extended_lut = "off";
defparam \src_data[14] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[14] .shared_arith = "off";

cyclonev_lcell_comb \src_data[22] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_22),
	.datad(!q_a_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22] .extended_lut = "off";
defparam \src_data[22] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[22] .shared_arith = "off";

cyclonev_lcell_comb \src_data[30] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_30),
	.datae(!q_a_30),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30] .extended_lut = "off";
defparam \src_data[30] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[30] .shared_arith = "off";

cyclonev_lcell_comb \src_data[5] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_5),
	.datae(!q_a_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5] .extended_lut = "off";
defparam \src_data[5] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[5] .shared_arith = "off";

cyclonev_lcell_comb \src_data[21] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_21),
	.datae(!q_a_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21] .extended_lut = "off";
defparam \src_data[21] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[21] .shared_arith = "off";

cyclonev_lcell_comb \src_data[4] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_4),
	.datad(!q_a_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4] .extended_lut = "off";
defparam \src_data[4] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[4] .shared_arith = "off";

cyclonev_lcell_comb \src_data[20] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_20),
	.datad(!q_a_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20] .extended_lut = "off";
defparam \src_data[20] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[20] .shared_arith = "off";

cyclonev_lcell_comb \src_data[3] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_3),
	.datae(!q_a_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3] .extended_lut = "off";
defparam \src_data[3] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[3] .shared_arith = "off";

cyclonev_lcell_comb \src_data[19] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_19),
	.datae(!q_a_19),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19] .extended_lut = "off";
defparam \src_data[19] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[19] .shared_arith = "off";

cyclonev_lcell_comb \src_data[1] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_1),
	.datad(!q_a_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1] .extended_lut = "off";
defparam \src_data[1] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[1] .shared_arith = "off";

cyclonev_lcell_comb \src_data[17] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!av_readdata_pre_17),
	.datad(!q_a_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17] .extended_lut = "off";
defparam \src_data[17] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[17] .shared_arith = "off";

cyclonev_lcell_comb \src_data[0] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_0),
	.datae(!q_a_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0] .extended_lut = "off";
defparam \src_data[0] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[16] (
	.dataa(!src0_valid),
	.datab(!src0_valid1),
	.datac(!\src_payload~0_combout ),
	.datad(!av_readdata_pre_16),
	.datae(!q_a_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16] .extended_lut = "off";
defparam \src_data[16] .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \src_data[16] .shared_arith = "off";

cyclonev_lcell_comb \src_payload~0 (
	.dataa(!hold_waitrequest),
	.datab(!read_latency_shift_reg_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\src_payload~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_payload~0 .extended_lut = "off";
defparam \src_payload~0 .lut_mask = 64'h7777777777777777;
defparam \src_payload~0 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_mm_interconnect_0_rsp_mux_001 (
	q_a_2,
	q_a_10,
	q_a_18,
	q_a_26,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_29,
	q_a_13,
	q_a_28,
	q_a_12,
	q_a_27,
	q_a_11,
	q_a_25,
	q_a_9,
	q_a_24,
	q_a_8,
	q_a_6,
	q_a_14,
	q_a_22,
	q_a_30,
	q_a_5,
	q_a_21,
	q_a_4,
	q_a_20,
	q_a_3,
	q_a_19,
	q_a_1,
	q_a_17,
	q_a_0,
	q_a_16,
	src1_valid,
	src1_valid1,
	WideOr11,
	av_readdata_pre_2,
	av_readdata_pre_10,
	av_readdata_pre_18,
	av_readdata_pre_26,
	av_readdata_pre_7,
	av_readdata_pre_23,
	av_readdata_pre_15,
	av_readdata_pre_31,
	av_readdata_pre_29,
	av_readdata_pre_13,
	av_readdata_pre_28,
	av_readdata_pre_12,
	av_readdata_pre_27,
	av_readdata_pre_11,
	av_readdata_pre_25,
	av_readdata_pre_9,
	av_readdata_pre_24,
	av_readdata_pre_8,
	av_readdata_pre_6,
	av_readdata_pre_14,
	av_readdata_pre_22,
	av_readdata_pre_30,
	av_readdata_pre_5,
	av_readdata_pre_21,
	av_readdata_pre_4,
	av_readdata_pre_20,
	av_readdata_pre_3,
	av_readdata_pre_19,
	av_readdata_pre_1,
	av_readdata_pre_17,
	av_readdata_pre_0,
	av_readdata_pre_16,
	src_data_5,
	src_data_3,
	src_data_1,
	src_data_4,
	src_data_2,
	src_data_28,
	src_data_31,
	src_data_27,
	src_data_29,
	src_data_30,
	src_data_0,
	src_data_23,
	src_data_26,
	src_data_22,
	src_data_24,
	src_data_25,
	src_data_16,
	src_data_15,
	src_data_13,
	src_data_14,
	src_data_12,
	src_data_11,
	src_data_8,
	src_data_19,
	src_data_18,
	src_data_17,
	src_data_10,
	src_data_9,
	src_data_21,
	src_data_20,
	src_data_7,
	src_data_6)/* synthesis synthesis_greybox=1 */;
input 	q_a_2;
input 	q_a_10;
input 	q_a_18;
input 	q_a_26;
input 	q_a_7;
input 	q_a_23;
input 	q_a_15;
input 	q_a_31;
input 	q_a_29;
input 	q_a_13;
input 	q_a_28;
input 	q_a_12;
input 	q_a_27;
input 	q_a_11;
input 	q_a_25;
input 	q_a_9;
input 	q_a_24;
input 	q_a_8;
input 	q_a_6;
input 	q_a_14;
input 	q_a_22;
input 	q_a_30;
input 	q_a_5;
input 	q_a_21;
input 	q_a_4;
input 	q_a_20;
input 	q_a_3;
input 	q_a_19;
input 	q_a_1;
input 	q_a_17;
input 	q_a_0;
input 	q_a_16;
input 	src1_valid;
input 	src1_valid1;
output 	WideOr11;
input 	av_readdata_pre_2;
input 	av_readdata_pre_10;
input 	av_readdata_pre_18;
input 	av_readdata_pre_26;
input 	av_readdata_pre_7;
input 	av_readdata_pre_23;
input 	av_readdata_pre_15;
input 	av_readdata_pre_31;
input 	av_readdata_pre_29;
input 	av_readdata_pre_13;
input 	av_readdata_pre_28;
input 	av_readdata_pre_12;
input 	av_readdata_pre_27;
input 	av_readdata_pre_11;
input 	av_readdata_pre_25;
input 	av_readdata_pre_9;
input 	av_readdata_pre_24;
input 	av_readdata_pre_8;
input 	av_readdata_pre_6;
input 	av_readdata_pre_14;
input 	av_readdata_pre_22;
input 	av_readdata_pre_30;
input 	av_readdata_pre_5;
input 	av_readdata_pre_21;
input 	av_readdata_pre_4;
input 	av_readdata_pre_20;
input 	av_readdata_pre_3;
input 	av_readdata_pre_19;
input 	av_readdata_pre_1;
input 	av_readdata_pre_17;
input 	av_readdata_pre_0;
input 	av_readdata_pre_16;
output 	src_data_5;
output 	src_data_3;
output 	src_data_1;
output 	src_data_4;
output 	src_data_2;
output 	src_data_28;
output 	src_data_31;
output 	src_data_27;
output 	src_data_29;
output 	src_data_30;
output 	src_data_0;
output 	src_data_23;
output 	src_data_26;
output 	src_data_22;
output 	src_data_24;
output 	src_data_25;
output 	src_data_16;
output 	src_data_15;
output 	src_data_13;
output 	src_data_14;
output 	src_data_12;
output 	src_data_11;
output 	src_data_8;
output 	src_data_19;
output 	src_data_18;
output 	src_data_17;
output 	src_data_10;
output 	src_data_9;
output 	src_data_21;
output 	src_data_20;
output 	src_data_7;
output 	src_data_6;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb WideOr1(
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(WideOr11),
	.sumout(),
	.cout(),
	.shareout());
defparam WideOr1.extended_lut = "off";
defparam WideOr1.lut_mask = 64'h7777777777777777;
defparam WideOr1.shared_arith = "off";

cyclonev_lcell_comb \src_data[5] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_5),
	.datad(!q_a_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_5),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[5] .extended_lut = "off";
defparam \src_data[5] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[5] .shared_arith = "off";

cyclonev_lcell_comb \src_data[3] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_3),
	.datad(!q_a_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_3),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[3] .extended_lut = "off";
defparam \src_data[3] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[3] .shared_arith = "off";

cyclonev_lcell_comb \src_data[1] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_1),
	.datad(!q_a_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_1),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[1] .extended_lut = "off";
defparam \src_data[1] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[1] .shared_arith = "off";

cyclonev_lcell_comb \src_data[4] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_4),
	.datad(!q_a_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_4),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[4] .extended_lut = "off";
defparam \src_data[4] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[4] .shared_arith = "off";

cyclonev_lcell_comb \src_data[2] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_2),
	.datad(!q_a_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_2),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[2] .extended_lut = "off";
defparam \src_data[2] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[2] .shared_arith = "off";

cyclonev_lcell_comb \src_data[28] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_28),
	.datad(!q_a_28),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_28),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[28] .extended_lut = "off";
defparam \src_data[28] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[28] .shared_arith = "off";

cyclonev_lcell_comb \src_data[31] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_31),
	.datad(!q_a_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_31),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[31] .extended_lut = "off";
defparam \src_data[31] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[31] .shared_arith = "off";

cyclonev_lcell_comb \src_data[27] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_27),
	.datad(!q_a_27),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_27),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[27] .extended_lut = "off";
defparam \src_data[27] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[27] .shared_arith = "off";

cyclonev_lcell_comb \src_data[29] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_29),
	.datad(!q_a_29),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_29),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[29] .extended_lut = "off";
defparam \src_data[29] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[29] .shared_arith = "off";

cyclonev_lcell_comb \src_data[30] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_30),
	.datad(!q_a_30),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_30),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[30] .extended_lut = "off";
defparam \src_data[30] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[30] .shared_arith = "off";

cyclonev_lcell_comb \src_data[0] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_0),
	.datad(!q_a_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_0),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[0] .extended_lut = "off";
defparam \src_data[0] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[0] .shared_arith = "off";

cyclonev_lcell_comb \src_data[23] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_23),
	.datad(!q_a_23),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_23),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[23] .extended_lut = "off";
defparam \src_data[23] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[23] .shared_arith = "off";

cyclonev_lcell_comb \src_data[26] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_26),
	.datad(!q_a_26),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_26),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[26] .extended_lut = "off";
defparam \src_data[26] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[26] .shared_arith = "off";

cyclonev_lcell_comb \src_data[22] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_22),
	.datad(!q_a_22),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_22),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[22] .extended_lut = "off";
defparam \src_data[22] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[22] .shared_arith = "off";

cyclonev_lcell_comb \src_data[24] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_24),
	.datad(!q_a_24),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_24),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[24] .extended_lut = "off";
defparam \src_data[24] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[24] .shared_arith = "off";

cyclonev_lcell_comb \src_data[25] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_25),
	.datad(!q_a_25),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_25),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[25] .extended_lut = "off";
defparam \src_data[25] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[25] .shared_arith = "off";

cyclonev_lcell_comb \src_data[16] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_16),
	.datad(!q_a_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_16),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[16] .extended_lut = "off";
defparam \src_data[16] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[16] .shared_arith = "off";

cyclonev_lcell_comb \src_data[15] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_15),
	.datad(!q_a_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_15),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[15] .extended_lut = "off";
defparam \src_data[15] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[15] .shared_arith = "off";

cyclonev_lcell_comb \src_data[13] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_13),
	.datad(!q_a_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_13),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[13] .extended_lut = "off";
defparam \src_data[13] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[13] .shared_arith = "off";

cyclonev_lcell_comb \src_data[14] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_14),
	.datad(!q_a_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_14),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[14] .extended_lut = "off";
defparam \src_data[14] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[14] .shared_arith = "off";

cyclonev_lcell_comb \src_data[12] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_12),
	.datad(!q_a_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_12),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[12] .extended_lut = "off";
defparam \src_data[12] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[12] .shared_arith = "off";

cyclonev_lcell_comb \src_data[11] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_11),
	.datad(!q_a_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_11),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[11] .extended_lut = "off";
defparam \src_data[11] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[11] .shared_arith = "off";

cyclonev_lcell_comb \src_data[8] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_8),
	.datad(!q_a_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_8),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[8] .extended_lut = "off";
defparam \src_data[8] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[8] .shared_arith = "off";

cyclonev_lcell_comb \src_data[19] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_19),
	.datad(!q_a_19),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_19),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[19] .extended_lut = "off";
defparam \src_data[19] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[19] .shared_arith = "off";

cyclonev_lcell_comb \src_data[18] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_18),
	.datad(!q_a_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_18),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[18] .extended_lut = "off";
defparam \src_data[18] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[18] .shared_arith = "off";

cyclonev_lcell_comb \src_data[17] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_17),
	.datad(!q_a_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_17),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[17] .extended_lut = "off";
defparam \src_data[17] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[17] .shared_arith = "off";

cyclonev_lcell_comb \src_data[10] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_10),
	.datad(!q_a_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_10),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[10] .extended_lut = "off";
defparam \src_data[10] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[10] .shared_arith = "off";

cyclonev_lcell_comb \src_data[9] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_9),
	.datad(!q_a_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_9),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[9] .extended_lut = "off";
defparam \src_data[9] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[9] .shared_arith = "off";

cyclonev_lcell_comb \src_data[21] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_21),
	.datad(!q_a_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_21),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[21] .extended_lut = "off";
defparam \src_data[21] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[21] .shared_arith = "off";

cyclonev_lcell_comb \src_data[20] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_20),
	.datad(!q_a_20),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_20),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[20] .extended_lut = "off";
defparam \src_data[20] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[20] .shared_arith = "off";

cyclonev_lcell_comb \src_data[7] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_7),
	.datad(!q_a_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_7),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[7] .extended_lut = "off";
defparam \src_data[7] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[7] .shared_arith = "off";

cyclonev_lcell_comb \src_data[6] (
	.dataa(!src1_valid),
	.datab(!src1_valid1),
	.datac(!av_readdata_pre_6),
	.datad(!q_a_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(src_data_6),
	.sumout(),
	.cout(),
	.shareout());
defparam \src_data[6] .extended_lut = "off";
defparam \src_data[6] .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \src_data[6] .shared_arith = "off";

endmodule

module embedded_system_embedded_system_nios2_qsys_0 (
	readdata_2,
	readdata_10,
	readdata_18,
	readdata_26,
	readdata_7,
	readdata_23,
	readdata_15,
	readdata_31,
	readdata_29,
	readdata_13,
	readdata_28,
	readdata_12,
	readdata_27,
	readdata_11,
	readdata_25,
	readdata_9,
	readdata_24,
	readdata_8,
	readdata_6,
	readdata_14,
	readdata_22,
	readdata_30,
	readdata_5,
	readdata_21,
	readdata_4,
	readdata_20,
	readdata_3,
	readdata_19,
	readdata_1,
	readdata_17,
	readdata_0,
	readdata_16,
	sr_0,
	ir_out_0,
	ir_out_1,
	r_sync_rst,
	hold_waitrequest,
	d_address_offset_field_0,
	d_write,
	d_address_tag_field_2,
	d_address_tag_field_1,
	d_address_tag_field_0,
	d_address_line_field_5,
	d_address_line_field_4,
	d_address_line_field_3,
	d_address_line_field_2,
	d_address_line_field_1,
	d_address_line_field_0,
	d_address_offset_field_2,
	d_address_offset_field_1,
	d_writedata_11,
	d_byteenable_0,
	d_writedata_10,
	d_writedata_9,
	d_writedata_8,
	d_writedata_13,
	d_writedata_12,
	d_writedata_21,
	d_writedata_20,
	d_writedata_25,
	d_writedata_17,
	d_writedata_24,
	d_writedata_16,
	d_writedata_27,
	d_writedata_19,
	d_writedata_26,
	d_writedata_18,
	d_writedata_23,
	d_writedata_15,
	d_writedata_22,
	d_writedata_14,
	d_read,
	suppress_change_dest_id,
	saved_grant_0,
	jtag_debug_module_waitrequest,
	mem_used_1,
	WideOr0,
	av_waitrequest,
	d_byteenable_1,
	d_writedata_2,
	d_writedata_0,
	d_writedata_3,
	d_writedata_1,
	hbreak_enabled1,
	i_read,
	src0_valid,
	ic_fill_tag_1,
	ic_fill_tag_0,
	ic_fill_line_6,
	Equal1,
	src0_valid1,
	src1_valid,
	saved_grant_1,
	rf_source_valid,
	d_writedata_6,
	d_writedata_4,
	d_writedata_7,
	d_writedata_5,
	r_early_rst,
	d_readdatavalid,
	suppress_change_dest_id1,
	WideOr01,
	WideOr02,
	nonposted_cmd_accepted,
	ic_fill_line_5,
	src_data_46,
	src_payload,
	ic_fill_ap_offset_0,
	src_data_38,
	ic_fill_line_1,
	src_data_42,
	ic_fill_line_0,
	src_data_41,
	ic_fill_ap_offset_2,
	src_data_40,
	ic_fill_ap_offset_1,
	src_data_39,
	ic_fill_line_4,
	src_data_45,
	ic_fill_line_3,
	src_data_44,
	ic_fill_line_2,
	src_data_43,
	src_payload1,
	src_data_32,
	src_payload2,
	src_payload3,
	WideOr1,
	d_readdata,
	jtag_debug_module_resetrequest,
	src_payload4,
	i_readdata,
	d_byteenable_2,
	d_byteenable_3,
	d_writedata_31,
	d_writedata_29,
	d_writedata_28,
	d_writedata_30,
	src_payload5,
	src_data_35,
	src_payload6,
	src_payload7,
	src_data_34,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_data_33,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	src_payload32,
	altera_internal_jtag,
	altera_internal_jtag1,
	NJQG9082,
	state_1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	irf_reg_1_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_2;
output 	readdata_10;
output 	readdata_18;
output 	readdata_26;
output 	readdata_7;
output 	readdata_23;
output 	readdata_15;
output 	readdata_31;
output 	readdata_29;
output 	readdata_13;
output 	readdata_28;
output 	readdata_12;
output 	readdata_27;
output 	readdata_11;
output 	readdata_25;
output 	readdata_9;
output 	readdata_24;
output 	readdata_8;
output 	readdata_6;
output 	readdata_14;
output 	readdata_22;
output 	readdata_30;
output 	readdata_5;
output 	readdata_21;
output 	readdata_4;
output 	readdata_20;
output 	readdata_3;
output 	readdata_19;
output 	readdata_1;
output 	readdata_17;
output 	readdata_0;
output 	readdata_16;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	r_sync_rst;
input 	hold_waitrequest;
output 	d_address_offset_field_0;
output 	d_write;
output 	d_address_tag_field_2;
output 	d_address_tag_field_1;
output 	d_address_tag_field_0;
output 	d_address_line_field_5;
output 	d_address_line_field_4;
output 	d_address_line_field_3;
output 	d_address_line_field_2;
output 	d_address_line_field_1;
output 	d_address_line_field_0;
output 	d_address_offset_field_2;
output 	d_address_offset_field_1;
output 	d_writedata_11;
output 	d_byteenable_0;
output 	d_writedata_10;
output 	d_writedata_9;
output 	d_writedata_8;
output 	d_writedata_13;
output 	d_writedata_12;
output 	d_writedata_21;
output 	d_writedata_20;
output 	d_writedata_25;
output 	d_writedata_17;
output 	d_writedata_24;
output 	d_writedata_16;
output 	d_writedata_27;
output 	d_writedata_19;
output 	d_writedata_26;
output 	d_writedata_18;
output 	d_writedata_23;
output 	d_writedata_15;
output 	d_writedata_22;
output 	d_writedata_14;
output 	d_read;
input 	suppress_change_dest_id;
input 	saved_grant_0;
output 	jtag_debug_module_waitrequest;
input 	mem_used_1;
input 	WideOr0;
input 	av_waitrequest;
output 	d_byteenable_1;
output 	d_writedata_2;
output 	d_writedata_0;
output 	d_writedata_3;
output 	d_writedata_1;
output 	hbreak_enabled1;
output 	i_read;
input 	src0_valid;
output 	ic_fill_tag_1;
output 	ic_fill_tag_0;
output 	ic_fill_line_6;
input 	Equal1;
input 	src0_valid1;
input 	src1_valid;
input 	saved_grant_1;
input 	rf_source_valid;
output 	d_writedata_6;
output 	d_writedata_4;
output 	d_writedata_7;
output 	d_writedata_5;
input 	r_early_rst;
input 	d_readdatavalid;
input 	suppress_change_dest_id1;
input 	WideOr01;
input 	WideOr02;
input 	nonposted_cmd_accepted;
output 	ic_fill_line_5;
input 	src_data_46;
input 	src_payload;
output 	ic_fill_ap_offset_0;
input 	src_data_38;
output 	ic_fill_line_1;
input 	src_data_42;
output 	ic_fill_line_0;
input 	src_data_41;
output 	ic_fill_ap_offset_2;
input 	src_data_40;
output 	ic_fill_ap_offset_1;
input 	src_data_39;
output 	ic_fill_line_4;
input 	src_data_45;
output 	ic_fill_line_3;
input 	src_data_44;
output 	ic_fill_line_2;
input 	src_data_43;
input 	src_payload1;
input 	src_data_32;
input 	src_payload2;
input 	src_payload3;
input 	WideOr1;
input 	[31:0] d_readdata;
output 	jtag_debug_module_resetrequest;
input 	src_payload4;
input 	[31:0] i_readdata;
output 	d_byteenable_2;
output 	d_byteenable_3;
output 	d_writedata_31;
output 	d_writedata_29;
output 	d_writedata_28;
output 	d_writedata_30;
input 	src_payload5;
input 	src_data_35;
input 	src_payload6;
input 	src_payload7;
input 	src_data_34;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_data_33;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	src_payload32;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	NJQG9082;
input 	state_1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[11] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[10] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[9] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[8] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[13] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[12] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[21] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[20] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[25] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[17] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[24] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[16] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[27] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[19] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[26] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[18] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[23] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[15] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[22] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[14] ;
wire \embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[1] ;
wire \embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[2] ;
wire \embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[3] ;
wire \embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[0] ;
wire \A_dc_xfer_wr_data[11]~q ;
wire \A_dc_xfer_wr_data[10]~q ;
wire \A_dc_xfer_wr_data[9]~q ;
wire \A_dc_xfer_wr_data[8]~q ;
wire \A_dc_xfer_wr_data[13]~q ;
wire \A_dc_xfer_wr_data[12]~q ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[2] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[0] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[3] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[1] ;
wire \A_dc_xfer_wr_data[21]~q ;
wire \A_dc_xfer_wr_data[20]~q ;
wire \A_dc_xfer_wr_data[25]~q ;
wire \A_dc_xfer_wr_data[17]~q ;
wire \A_dc_xfer_wr_data[24]~q ;
wire \A_dc_xfer_wr_data[16]~q ;
wire \A_dc_xfer_wr_data[27]~q ;
wire \A_dc_xfer_wr_data[19]~q ;
wire \A_dc_xfer_wr_data[26]~q ;
wire \A_dc_xfer_wr_data[18]~q ;
wire \A_dc_xfer_wr_data[23]~q ;
wire \A_dc_xfer_wr_data[15]~q ;
wire \A_dc_xfer_wr_data[22]~q ;
wire \A_dc_xfer_wr_data[14]~q ;
wire \embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[4] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[2] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[2] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[13] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[13] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[12] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[12] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[11] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[11] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[10] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[10] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[9] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[9] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[8] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[8] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[7] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[7] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[6] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[6] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[5] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[5] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[4] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[4] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[3] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[3] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[1] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[0] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ;
wire \A_dc_xfer_wr_data[2]~q ;
wire \A_dc_xfer_wr_data[0]~q ;
wire \A_dc_xfer_wr_data[3]~q ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[6] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[4] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[7] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[5] ;
wire \A_dc_xfer_wr_data[1]~q ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[21] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[20] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[25] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[17] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[24] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[16] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[27] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[19] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[26] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[18] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[23] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[15] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[22] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[14] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[5] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[3] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[4] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ;
wire \embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[0] ;
wire \embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[1] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[27] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[29] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[29] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[30] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[30] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[31] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[31] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[17] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[16] ;
wire \embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[28] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[28] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[18] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[26] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[19] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[21] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[15] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[25] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[20] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[22] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[14] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[24] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[23] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[1] ;
wire \embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[0] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[16] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[15] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[13] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[14] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[8] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ;
wire \embedded_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[1] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[19] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[18] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[17] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[10] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[9] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ;
wire \embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ;
wire \A_dc_xfer_wr_data[6]~q ;
wire \A_dc_xfer_wr_data[4]~q ;
wire \A_dc_xfer_wr_data[7]~q ;
wire \A_dc_xfer_wr_data[5]~q ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[21] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[20] ;
wire \embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[7] ;
wire \embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[9] ;
wire \embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[6] ;
wire \embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[8] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[7] ;
wire \embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[6] ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~1_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~5_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~9_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~13_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~17_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~21_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~25_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~29_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~33_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~37_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~41_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~45_sumout ;
wire \ic_fill_valid_bits[5]~q ;
wire \ic_fill_valid_bits[7]~q ;
wire \ic_fill_valid_bits[4]~q ;
wire \embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[3] ;
wire \embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[5] ;
wire \embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[2] ;
wire \embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[4] ;
wire \ic_fill_valid_bits[6]~q ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~49_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~53_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~57_sumout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|Add0~61_sumout ;
wire \ic_fill_valid_bits[1]~q ;
wire \ic_fill_valid_bits[3]~q ;
wire \ic_fill_valid_bits[0]~q ;
wire \ic_fill_valid_bits[2]~q ;
wire \A_mul_src2[0]~q ;
wire \A_mul_src2[1]~q ;
wire \A_mul_src2[2]~q ;
wire \A_mul_src2[3]~q ;
wire \A_mul_src2[4]~q ;
wire \A_mul_src2[5]~q ;
wire \A_mul_src2[6]~q ;
wire \A_mul_src2[7]~q ;
wire \A_mul_src2[8]~q ;
wire \A_mul_src2[9]~q ;
wire \A_mul_src2[10]~q ;
wire \A_mul_src2[11]~q ;
wire \A_mul_src2[12]~q ;
wire \A_mul_src2[13]~q ;
wire \A_mul_src2[14]~q ;
wire \A_mul_src2[15]~q ;
wire \A_mul_src1[0]~q ;
wire \A_mul_src1[1]~q ;
wire \A_mul_src1[2]~q ;
wire \A_mul_src1[3]~q ;
wire \A_mul_src1[4]~q ;
wire \A_mul_src1[5]~q ;
wire \A_mul_src1[6]~q ;
wire \A_mul_src1[7]~q ;
wire \A_mul_src1[8]~q ;
wire \A_mul_src1[9]~q ;
wire \A_mul_src1[10]~q ;
wire \A_mul_src1[11]~q ;
wire \A_mul_src1[12]~q ;
wire \A_mul_src1[13]~q ;
wire \A_mul_src1[14]~q ;
wire \A_mul_src1[15]~q ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[31] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[29] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[28] ;
wire \embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[30] ;
wire \A_mul_src2[16]~q ;
wire \A_mul_src2[17]~q ;
wire \A_mul_src2[18]~q ;
wire \A_mul_src2[19]~q ;
wire \A_mul_src2[20]~q ;
wire \A_mul_src2[21]~q ;
wire \A_mul_src2[22]~q ;
wire \A_mul_src2[23]~q ;
wire \A_mul_src2[24]~q ;
wire \A_mul_src2[25]~q ;
wire \A_mul_src2[26]~q ;
wire \A_mul_src2[27]~q ;
wire \A_mul_src2[28]~q ;
wire \A_mul_src2[29]~q ;
wire \A_mul_src2[30]~q ;
wire \A_mul_src2[31]~q ;
wire \embedded_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[0] ;
wire \A_dc_xfer_wr_data[31]~q ;
wire \A_dc_xfer_wr_data[29]~q ;
wire \A_dc_xfer_wr_data[28]~q ;
wire \A_dc_xfer_wr_data[30]~q ;
wire \A_mul_src1[16]~q ;
wire \A_mul_src1[17]~q ;
wire \A_mul_src1[18]~q ;
wire \A_mul_src1[19]~q ;
wire \A_mul_src1[20]~q ;
wire \A_mul_src1[21]~q ;
wire \A_mul_src1[22]~q ;
wire \A_mul_src1[23]~q ;
wire \A_mul_src1[24]~q ;
wire \A_mul_src1[25]~q ;
wire \A_mul_src1[26]~q ;
wire \A_mul_src1[27]~q ;
wire \A_mul_src1[28]~q ;
wire \A_mul_src1[29]~q ;
wire \A_mul_src1[30]~q ;
wire \A_mul_src1[31]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_oci_debug|jtag_break~q ;
wire \A_dc_xfer_wr_active~q ;
wire \A_dc_wb_rd_en~0_combout ;
wire \A_dc_wb_rd_en~combout ;
wire \A_dc_xfer_wr_offset[0]~q ;
wire \A_dc_xfer_wr_offset[1]~q ;
wire \A_dc_xfer_wr_offset[2]~q ;
wire \A_dc_wb_rd_addr_offset[0]~q ;
wire \A_dc_wb_rd_addr_offset[1]~q ;
wire \A_dc_wb_rd_addr_offset[2]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_single_step_mode~q ;
wire \A_dc_fill_starting_d1~q ;
wire \A_en_d1~q ;
wire \A_ctrl_dc_index_inv~q ;
wire \A_ctrl_dc_addr_inv~q ;
wire \dc_tag_wr_port_addr~0_combout ;
wire \dc_tag_wr_port_en~combout ;
wire \dc_tag_wr_port_data[1]~0_combout ;
wire \dc_tag_wr_port_addr[0]~1_combout ;
wire \dc_tag_wr_port_addr[1]~2_combout ;
wire \dc_tag_wr_port_addr[2]~3_combout ;
wire \dc_tag_wr_port_addr[3]~4_combout ;
wire \dc_tag_wr_port_addr[4]~5_combout ;
wire \dc_tag_wr_port_addr[5]~6_combout ;
wire \dc_tag_rd_port_addr[0]~0_combout ;
wire \dc_tag_rd_port_addr[1]~1_combout ;
wire \dc_tag_rd_port_addr[2]~2_combout ;
wire \dc_tag_rd_port_addr[3]~3_combout ;
wire \dc_tag_rd_port_addr[4]~4_combout ;
wire \dc_tag_rd_port_addr[5]~5_combout ;
wire \dc_tag_wr_port_data[2]~1_combout ;
wire \dc_tag_wr_port_data[3]~2_combout ;
wire \dc_tag_wr_port_data[0]~3_combout ;
wire \A_dc_xfer_rd_data_active~q ;
wire \A_dc_rd_data[11]~q ;
wire \A_dc_xfer_rd_data_offset_match~q ;
wire \A_dc_xfer_wr_offset_nxt[0]~0_combout ;
wire \A_dc_xfer_wr_offset_nxt[1]~1_combout ;
wire \A_dc_xfer_wr_offset_nxt[2]~2_combout ;
wire \A_dc_wb_rd_addr_offset_nxt[0]~0_combout ;
wire \A_dc_wb_rd_addr_offset_nxt[1]~1_combout ;
wire \A_dc_wb_rd_addr_offset_nxt[2]~2_combout ;
wire \A_dc_rd_data[10]~q ;
wire \A_dc_rd_data[9]~q ;
wire \A_dc_rd_data[8]~q ;
wire \A_dc_rd_data[13]~q ;
wire \A_dc_rd_data[12]~q ;
wire \A_dc_rd_data[21]~q ;
wire \A_dc_rd_data[20]~q ;
wire \A_dc_rd_data[25]~q ;
wire \A_dc_rd_data[17]~q ;
wire \A_dc_rd_data[24]~q ;
wire \A_dc_rd_data[16]~q ;
wire \A_dc_rd_data[27]~q ;
wire \A_dc_rd_data[19]~q ;
wire \A_dc_rd_data[26]~q ;
wire \A_dc_rd_data[18]~q ;
wire \A_dc_rd_data[23]~q ;
wire \A_dc_rd_data[15]~q ;
wire \A_dc_rd_data[22]~q ;
wire \A_dc_rd_data[14]~q ;
wire \M_ctrl_dc_index_inv~q ;
wire \M_ctrl_dc_addr_inv~q ;
wire \A_valid_st_writes_mem~q ;
wire \dc_tag_wr_port_data[4]~4_combout ;
wire \rf_b_rd_port_addr[0]~0_combout ;
wire \rf_b_rd_port_addr[1]~1_combout ;
wire \rf_b_rd_port_addr[2]~2_combout ;
wire \rf_b_rd_port_addr[3]~3_combout ;
wire \rf_b_rd_port_addr[4]~4_combout ;
wire \rf_a_rd_port_addr[0]~0_combout ;
wire \rf_a_rd_port_addr[1]~1_combout ;
wire \rf_a_rd_port_addr[2]~2_combout ;
wire \rf_a_rd_port_addr[3]~3_combout ;
wire \rf_a_rd_port_addr[4]~4_combout ;
wire \A_dc_valid_st_bypass_hit_wr_en~combout ;
wire \dc_data_wr_port_en~combout ;
wire \M_dc_st_data[11]~0_combout ;
wire \A_dc_st_data[11]~q ;
wire \A_ctrl_st~q ;
wire \dc_data_wr_port_data[13]~0_combout ;
wire \dc_data_wr_port_data[11]~1_combout ;
wire \dc_data_wr_port_addr[0]~0_combout ;
wire \dc_data_wr_port_addr[1]~1_combout ;
wire \dc_data_wr_port_addr[2]~2_combout ;
wire \dc_data_wr_port_addr[3]~3_combout ;
wire \dc_data_wr_port_addr[4]~4_combout ;
wire \dc_data_wr_port_addr[5]~5_combout ;
wire \dc_data_wr_port_addr[6]~6_combout ;
wire \dc_data_wr_port_addr[7]~7_combout ;
wire \dc_data_wr_port_addr[8]~8_combout ;
wire \dc_data_rd_port_addr[0]~0_combout ;
wire \dc_data_rd_port_addr[1]~1_combout ;
wire \dc_data_rd_port_addr[2]~2_combout ;
wire \dc_data_rd_port_addr[3]~3_combout ;
wire \dc_data_rd_port_addr[4]~4_combout ;
wire \dc_data_rd_port_addr[5]~5_combout ;
wire \dc_data_rd_port_addr[6]~6_combout ;
wire \dc_data_rd_port_addr[7]~7_combout ;
wire \dc_data_rd_port_addr[8]~8_combout ;
wire \A_dc_xfer_rd_addr_offset_match~0_combout ;
wire \A_dc_xfer_rd_addr_offset_match~combout ;
wire \M_dc_st_data[10]~1_combout ;
wire \A_dc_st_data[10]~q ;
wire \dc_data_wr_port_data[10]~2_combout ;
wire \M_dc_st_data[9]~2_combout ;
wire \A_dc_st_data[9]~q ;
wire \dc_data_wr_port_data[9]~3_combout ;
wire \M_dc_st_data[8]~3_combout ;
wire \A_dc_st_data[8]~q ;
wire \dc_data_wr_port_data[8]~4_combout ;
wire \M_dc_st_data[13]~4_combout ;
wire \A_dc_st_data[13]~q ;
wire \dc_data_wr_port_data[13]~5_combout ;
wire \M_dc_st_data[12]~5_combout ;
wire \A_dc_st_data[12]~q ;
wire \dc_data_wr_port_data[12]~6_combout ;
wire \A_dc_rd_data[2]~q ;
wire \A_dc_rd_data[0]~q ;
wire \A_dc_rd_data[3]~q ;
wire \A_dc_rd_data[1]~q ;
wire \M_dc_st_data[21]~6_combout ;
wire \A_dc_st_data[21]~q ;
wire \dc_data_wr_port_data[18]~7_combout ;
wire \dc_data_wr_port_data[21]~8_combout ;
wire \M_dc_st_data[20]~7_combout ;
wire \A_dc_st_data[20]~q ;
wire \dc_data_wr_port_data[20]~9_combout ;
wire \M_dc_st_data[25]~8_combout ;
wire \A_dc_st_data[25]~q ;
wire \dc_data_wr_port_data[25]~10_combout ;
wire \dc_data_wr_port_data[25]~11_combout ;
wire \M_dc_st_data[17]~9_combout ;
wire \A_dc_st_data[17]~q ;
wire \dc_data_wr_port_data[17]~12_combout ;
wire \M_dc_st_data[24]~10_combout ;
wire \A_dc_st_data[24]~q ;
wire \dc_data_wr_port_data[24]~13_combout ;
wire \M_dc_st_data[16]~11_combout ;
wire \A_dc_st_data[16]~q ;
wire \dc_data_wr_port_data[16]~14_combout ;
wire \M_dc_st_data[27]~12_combout ;
wire \A_dc_st_data[27]~q ;
wire \dc_data_wr_port_data[27]~15_combout ;
wire \M_dc_st_data[19]~13_combout ;
wire \A_dc_st_data[19]~q ;
wire \dc_data_wr_port_data[19]~16_combout ;
wire \M_dc_st_data[26]~14_combout ;
wire \A_dc_st_data[26]~q ;
wire \dc_data_wr_port_data[26]~17_combout ;
wire \M_dc_st_data[18]~15_combout ;
wire \A_dc_st_data[18]~q ;
wire \dc_data_wr_port_data[18]~18_combout ;
wire \M_dc_st_data[23]~16_combout ;
wire \A_dc_st_data[23]~q ;
wire \dc_data_wr_port_data[23]~19_combout ;
wire \M_dc_st_data[15]~17_combout ;
wire \A_dc_st_data[15]~q ;
wire \dc_data_wr_port_data[15]~20_combout ;
wire \M_dc_st_data[22]~18_combout ;
wire \A_dc_st_data[22]~q ;
wire \dc_data_wr_port_data[22]~21_combout ;
wire \M_dc_st_data[14]~19_combout ;
wire \A_dc_st_data[14]~q ;
wire \dc_data_wr_port_data[14]~22_combout ;
wire \i_readdata_d1[5]~q ;
wire \i_readdata_d1[3]~q ;
wire \i_readdata_d1[1]~q ;
wire \i_readdata_d1[4]~q ;
wire \i_readdata_d1[2]~q ;
wire \i_readdata_d1[28]~q ;
wire \i_readdata_d1[31]~q ;
wire \i_readdata_d1[27]~q ;
wire \i_readdata_d1[29]~q ;
wire \i_readdata_d1[30]~q ;
wire \i_readdata_d1[0]~q ;
wire \i_readdata_d1[23]~q ;
wire \i_readdata_d1[26]~q ;
wire \i_readdata_d1[22]~q ;
wire \i_readdata_d1[24]~q ;
wire \i_readdata_d1[25]~q ;
wire \ic_tag_clr_valid_bits~q ;
wire \ic_tag_wren~combout ;
wire \ic_tag_wraddress[0]~q ;
wire \ic_tag_wraddress[1]~q ;
wire \ic_tag_wraddress[2]~q ;
wire \ic_tag_wraddress[3]~q ;
wire \ic_tag_wraddress[4]~q ;
wire \ic_tag_wraddress[5]~q ;
wire \ic_tag_wraddress[6]~q ;
wire \i_readdata_d1[16]~q ;
wire \i_readdata_d1[15]~q ;
wire \i_readdata_d1[13]~q ;
wire \i_readdata_d1[14]~q ;
wire \i_readdata_d1[12]~q ;
wire \i_readdata_d1[11]~q ;
wire \E_ctrl_dc_index_inv~0_combout ;
wire \M_ctrl_st~q ;
wire \M_valid_st_writes_mem~combout ;
wire \i_readdata_d1[8]~q ;
wire \M_dc_st_data[2]~20_combout ;
wire \A_dc_st_data[2]~q ;
wire \dc_data_wr_port_data[1]~23_combout ;
wire \dc_data_wr_port_data[2]~24_combout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ;
wire \M_ctrl_br_cond~q ;
wire \M_bht_wr_en_unfiltered~combout ;
wire \M_bht_data[1]~q ;
wire \M_bht_data[0]~q ;
wire \M_br_mispredict~q ;
wire \M_bht_wr_data_unfiltered[1]~0_combout ;
wire \M_bht_ptr_unfiltered[0]~q ;
wire \M_bht_ptr_unfiltered[1]~q ;
wire \M_bht_ptr_unfiltered[2]~q ;
wire \M_bht_ptr_unfiltered[3]~q ;
wire \M_bht_ptr_unfiltered[4]~q ;
wire \M_bht_ptr_unfiltered[5]~q ;
wire \M_bht_ptr_unfiltered[6]~q ;
wire \M_bht_ptr_unfiltered[7]~q ;
wire \M_br_cond_taken_history[0]~q ;
wire \F_bht_ptr_nxt[0]~combout ;
wire \M_br_cond_taken_history[1]~q ;
wire \F_bht_ptr_nxt[1]~combout ;
wire \M_br_cond_taken_history[2]~q ;
wire \F_bht_ptr_nxt[2]~combout ;
wire \M_br_cond_taken_history[3]~q ;
wire \F_bht_ptr_nxt[3]~combout ;
wire \M_br_cond_taken_history[4]~q ;
wire \F_bht_ptr_nxt[4]~combout ;
wire \M_br_cond_taken_history[5]~q ;
wire \F_bht_ptr_nxt[5]~combout ;
wire \M_br_cond_taken_history[6]~q ;
wire \F_bht_ptr_nxt[6]~combout ;
wire \M_br_cond_taken_history[7]~q ;
wire \F_bht_ptr_nxt[7]~combout ;
wire \i_readdata_d1[19]~q ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ;
wire \M_dc_st_data[29]~21_combout ;
wire \A_dc_st_data[29]~q ;
wire \dc_data_wr_port_data[29]~25_combout ;
wire \M_dc_st_data[7]~22_combout ;
wire \A_dc_st_data[7]~q ;
wire \dc_data_wr_port_data[7]~26_combout ;
wire \M_dc_st_data[31]~23_combout ;
wire \A_dc_st_data[31]~q ;
wire \dc_data_wr_port_data[31]~27_combout ;
wire \i_readdata_d1[18]~q ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ;
wire \M_dc_st_data[28]~24_combout ;
wire \A_dc_st_data[28]~q ;
wire \dc_data_wr_port_data[28]~28_combout ;
wire \i_readdata_d1[17]~q ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ;
wire \M_dc_st_data[6]~25_combout ;
wire \A_dc_st_data[6]~q ;
wire \dc_data_wr_port_data[6]~29_combout ;
wire \M_dc_st_data[30]~26_combout ;
wire \A_dc_st_data[30]~q ;
wire \dc_data_wr_port_data[30]~30_combout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ;
wire \M_dc_st_data[5]~27_combout ;
wire \A_dc_st_data[5]~q ;
wire \dc_data_wr_port_data[5]~31_combout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ;
wire \i_readdata_d1[10]~q ;
wire \M_dc_st_data[4]~28_combout ;
wire \A_dc_st_data[4]~q ;
wire \dc_data_wr_port_data[4]~32_combout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ;
wire \i_readdata_d1[9]~q ;
wire \M_dc_st_data[3]~29_combout ;
wire \A_dc_st_data[3]~q ;
wire \dc_data_wr_port_data[3]~33_combout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ;
wire \M_dc_st_data[1]~30_combout ;
wire \A_dc_st_data[1]~q ;
wire \dc_data_wr_port_data[1]~34_combout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ;
wire \M_dc_st_data[0]~31_combout ;
wire \A_dc_st_data[0]~q ;
wire \dc_data_wr_port_data[0]~35_combout ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ;
wire \A_dc_rd_data[6]~q ;
wire \A_dc_rd_data[4]~q ;
wire \A_dc_rd_data[7]~q ;
wire \A_dc_rd_data[5]~q ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ;
wire \the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ;
wire \i_readdata_d1[21]~q ;
wire \i_readdata_d1[20]~q ;
wire \clr_break_line~q ;
wire \ic_tag_clr_valid_bits_nxt~combout ;
wire \ic_tag_wraddress_nxt~7_combout ;
wire \ic_tag_wraddress_nxt[0]~8_combout ;
wire \ic_tag_wraddress_nxt[1]~9_combout ;
wire \ic_tag_wraddress_nxt[1]~10_combout ;
wire \ic_tag_wraddress_nxt[2]~11_combout ;
wire \ic_tag_wraddress_nxt[3]~12_combout ;
wire \ic_tag_wraddress_nxt[4]~13_combout ;
wire \ic_tag_wraddress_nxt[5]~14_combout ;
wire \ic_tag_wraddress_nxt[6]~15_combout ;
wire \i_readdata_d1[7]~q ;
wire \i_readdata_d1[6]~q ;
wire \E_bht_data[0]~q ;
wire \E_br_mispredict~combout ;
wire \E_bht_ptr[0]~q ;
wire \E_bht_ptr[1]~q ;
wire \E_bht_ptr[2]~q ;
wire \E_bht_ptr[3]~q ;
wire \E_bht_ptr[4]~q ;
wire \E_bht_ptr[5]~q ;
wire \E_bht_ptr[6]~q ;
wire \E_bht_ptr[7]~q ;
wire \M_br_cond_taken_history[0]~0_combout ;
wire \M_br_cond_taken_history[0]~1_combout ;
wire \ic_fill_valid_bits_nxt~0_combout ;
wire \ic_fill_valid_bits_en~combout ;
wire \ic_fill_valid_bits_nxt~1_combout ;
wire \ic_fill_valid_bits_nxt~2_combout ;
wire \ic_fill_valid_bits_nxt~3_combout ;
wire \D_bht_data[0]~q ;
wire \D_bht_ptr[0]~q ;
wire \D_bht_ptr[1]~q ;
wire \D_bht_ptr[2]~q ;
wire \D_bht_ptr[3]~q ;
wire \D_bht_ptr[4]~q ;
wire \D_bht_ptr[5]~q ;
wire \D_bht_ptr[6]~q ;
wire \D_bht_ptr[7]~q ;
wire \ic_fill_valid_bits_nxt~4_combout ;
wire \ic_fill_valid_bits_nxt~5_combout ;
wire \ic_fill_valid_bits_nxt~6_combout ;
wire \ic_fill_valid_bits_nxt~7_combout ;
wire \M_src2[0]~q ;
wire \M_src2[1]~q ;
wire \M_src2[2]~q ;
wire \M_src2[3]~q ;
wire \M_src2[4]~q ;
wire \M_src2[5]~q ;
wire \M_src2[6]~q ;
wire \M_src2[7]~q ;
wire \M_src2[8]~q ;
wire \M_src2[9]~q ;
wire \M_src2[10]~q ;
wire \M_src2[11]~q ;
wire \M_src2[12]~q ;
wire \M_src2[13]~q ;
wire \M_src2[14]~q ;
wire \M_src2[15]~q ;
wire \M_src1[0]~q ;
wire \M_src1[1]~q ;
wire \M_src1[2]~q ;
wire \M_src1[3]~q ;
wire \M_src1[4]~q ;
wire \M_src1[5]~q ;
wire \M_src1[6]~q ;
wire \M_src1[7]~q ;
wire \M_src1[8]~q ;
wire \M_src1[9]~q ;
wire \M_src1[10]~q ;
wire \M_src1[11]~q ;
wire \M_src1[12]~q ;
wire \M_src1[13]~q ;
wire \M_src1[14]~q ;
wire \M_src1[15]~q ;
wire \F_bht_ptr[0]~q ;
wire \F_bht_ptr[1]~q ;
wire \F_bht_ptr[2]~q ;
wire \F_bht_ptr[3]~q ;
wire \F_bht_ptr[4]~q ;
wire \F_bht_ptr[5]~q ;
wire \F_bht_ptr[6]~q ;
wire \F_bht_ptr[7]~q ;
wire \M_src2[16]~q ;
wire \M_src2[17]~q ;
wire \M_src2[18]~q ;
wire \M_src2[19]~q ;
wire \M_src2[20]~q ;
wire \M_src2[21]~q ;
wire \M_src2[22]~q ;
wire \M_src2[23]~q ;
wire \M_src2[24]~q ;
wire \M_src2[25]~q ;
wire \M_src2[26]~q ;
wire \M_src2[27]~q ;
wire \M_src2[28]~q ;
wire \M_src2[29]~q ;
wire \M_src2[30]~q ;
wire \M_src2[31]~q ;
wire \A_dc_rd_data[31]~q ;
wire \A_dc_rd_data[29]~q ;
wire \A_dc_rd_data[28]~q ;
wire \A_dc_rd_data[30]~q ;
wire \M_src1[16]~q ;
wire \M_src1[17]~q ;
wire \M_src1[18]~q ;
wire \M_src1[19]~q ;
wire \M_src1[20]~q ;
wire \M_src1[21]~q ;
wire \M_src1[22]~q ;
wire \M_src1[23]~q ;
wire \M_src1[24]~q ;
wire \M_src1[25]~q ;
wire \M_src1[26]~q ;
wire \M_src1[27]~q ;
wire \M_src1[28]~q ;
wire \M_src1[29]~q ;
wire \M_src1[30]~q ;
wire \M_src1[31]~q ;
wire \ic_tag_clr_valid_bits~0_combout ;
wire \M_br_mispredict~_wirecell_combout ;
wire \A_dc_wb_wr_starting~combout ;
wire \av_wr_data_transfer~0_combout ;
wire \A_dc_wr_data_cnt_nxt[0]~3_combout ;
wire \hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ;
wire \A_dc_wb_wr_active_nxt~0_combout ;
wire \A_dc_wb_wr_active~q ;
wire \A_dc_wr_data_cnt[2]~0_combout ;
wire \A_dc_wr_data_cnt[0]~q ;
wire \A_dc_wr_data_cnt_nxt[1]~2_combout ;
wire \A_dc_wr_data_cnt[1]~q ;
wire \A_dc_wr_data_cnt_nxt[2]~1_combout ;
wire \A_dc_wr_data_cnt[2]~q ;
wire \A_dc_wr_data_cnt_nxt[3]~0_combout ;
wire \A_dc_wr_data_cnt[3]~q ;
wire \A_dc_wb_active_nxt~0_combout ;
wire \A_dc_wb_active~q ;
wire \E_iw[0]~q ;
wire \F_iw[5]~1_combout ;
wire \F_iw[3]~2_combout ;
wire \F_iw[1]~3_combout ;
wire \F_iw[4]~4_combout ;
wire \F_iw[2]~5_combout ;
wire \F_ctrl_a_not_src~0_combout ;
wire \D_ctrl_a_not_src~q ;
wire \F_ctrl_b_is_dst~0_combout ;
wire \D_ctrl_b_is_dst~q ;
wire \M_ctrl_late_result~q ;
wire \F_iw[19]~13_combout ;
wire \D_iw[19]~q ;
wire \D_iw[24]~q ;
wire \F_ctrl_implicit_dst_retaddr~0_combout ;
wire \D_ctrl_implicit_dst_retaddr~q ;
wire \F_iw[13]~8_combout ;
wire \F_ctrl_implicit_dst_eretaddr~0_combout ;
wire \Equal2~0_combout ;
wire \F_ctrl_implicit_dst_eretaddr~1_combout ;
wire \D_ctrl_implicit_dst_eretaddr~q ;
wire \D_dst_regnum[2]~3_combout ;
wire \E_dst_regnum[2]~q ;
wire \F_iw[16]~6_combout ;
wire \D_iw[16]~q ;
wire \E_iw[16]~q ;
wire \F_iw[15]~7_combout ;
wire \D_iw[15]~q ;
wire \E_iw[15]~q ;
wire \D_iw[13]~q ;
wire \E_iw[13]~q ;
wire \E_hbreak_req~0_combout ;
wire \D_iw[3]~q ;
wire \E_iw[3]~q ;
wire \D_iw[1]~q ;
wire \E_iw[1]~q ;
wire \D_iw[4]~q ;
wire \E_iw[4]~q ;
wire \D_iw[2]~q ;
wire \E_iw[2]~q ;
wire \Equal209~0_combout ;
wire \F_iw[14]~10_combout ;
wire \D_iw[14]~q ;
wire \E_iw[14]~q ;
wire \F_iw[12]~11_combout ;
wire \D_iw[12]~q ;
wire \E_iw[12]~q ;
wire \F_iw[11]~12_combout ;
wire \D_iw[11]~q ;
wire \E_iw[11]~q ;
wire \E_hbreak_req~1_combout ;
wire \E_hbreak_req~combout ;
wire \D_bht_data[1]~q ;
wire \E_bht_data[1]~q ;
wire \D_ctrl_cmp~3_combout ;
wire \D_ctrl_alu_subtract~0_combout ;
wire \D_ctrl_alu_subtract~1_combout ;
wire \D_ctrl_alu_subtract~2_combout ;
wire \E_ctrl_alu_subtract~q ;
wire \Equal154~1_combout ;
wire \Equal154~3_combout ;
wire \D_ctrl_alu_signed_comparison~0_combout ;
wire \D_ctrl_alu_signed_comparison~1_combout ;
wire \E_ctrl_alu_signed_comparison~q ;
wire \F_ctrl_src2_choose_imm~0_combout ;
wire \F_ctrl_src2_choose_imm~combout ;
wire \D_ctrl_src2_choose_imm~q ;
wire \D_iw[23]~q ;
wire \F_iw[18]~14_combout ;
wire \D_iw[18]~q ;
wire \D_dst_regnum[1]~0_combout ;
wire \D_iw[26]~q ;
wire \F_iw[21]~15_combout ;
wire \D_iw[21]~q ;
wire \D_dst_regnum[4]~1_combout ;
wire \F_ctrl_ignore_dst~combout ;
wire \D_ctrl_ignore_dst~q ;
wire \D_iw[22]~q ;
wire \D_iw[17]~q ;
wire \D_dst_regnum[0]~2_combout ;
wire \D_iw[25]~q ;
wire \F_iw[20]~16_combout ;
wire \D_iw[20]~q ;
wire \D_dst_regnum[3]~4_combout ;
wire \Equal295~0_combout ;
wire \D_wr_dst_reg~combout ;
wire \D_regnum_b_cmp_F~0_combout ;
wire \D_regnum_b_cmp_F~combout ;
wire \E_regnum_b_cmp_D~q ;
wire \E_dst_regnum[4]~q ;
wire \M_dst_regnum[4]~q ;
wire \M_wr_dst_reg_from_E~q ;
wire \E_dst_regnum[0]~q ;
wire \M_dst_regnum[0]~q ;
wire \E_dst_regnum[1]~q ;
wire \M_dst_regnum[1]~q ;
wire \M_regnum_b_cmp_F~0_combout ;
wire \M_dst_regnum[2]~q ;
wire \E_dst_regnum[3]~q ;
wire \M_dst_regnum[3]~q ;
wire \M_regnum_b_cmp_F~1_combout ;
wire \M_regnum_b_cmp_F~combout ;
wire \A_regnum_b_cmp_D~q ;
wire \A_dst_regnum_from_M[4]~q ;
wire \A_wr_dst_reg_from_M~q ;
wire \A_dst_regnum_from_M[0]~q ;
wire \A_dst_regnum_from_M[1]~q ;
wire \A_regnum_b_cmp_F~0_combout ;
wire \A_dst_regnum_from_M[2]~q ;
wire \A_dst_regnum_from_M[3]~q ;
wire \A_regnum_b_cmp_F~1_combout ;
wire \A_regnum_b_cmp_F~combout ;
wire \W_regnum_b_cmp_D~q ;
wire \D_src2_reg[5]~0_combout ;
wire \Equal297~0_combout ;
wire \D_src2_reg[5]~1_combout ;
wire \D_src2_reg[5]~2_combout ;
wire \D_src2_reg[0]~55_combout ;
wire \Equal92~0_combout ;
wire \D_ctrl_logic~0_combout ;
wire \D_ctrl_logic~1_combout ;
wire \D_ctrl_logic~2_combout ;
wire \E_ctrl_logic~q ;
wire \Equal105~0_combout ;
wire \Equal154~0_combout ;
wire \D_ctrl_retaddr~1_combout ;
wire \D_ctrl_retaddr~0_combout ;
wire \E_ctrl_retaddr~q ;
wire \D_ctrl_cmp~2_combout ;
wire \D_ctrl_cmp~0_combout ;
wire \D_ctrl_cmp~1_combout ;
wire \E_ctrl_cmp~q ;
wire \E_alu_result~0_combout ;
wire \D_ctrl_late_result~3_combout ;
wire \D_ctrl_mul_lsw~0_combout ;
wire \E_ctrl_mul_lsw~q ;
wire \M_ctrl_mul_lsw~q ;
wire \A_ctrl_mul_lsw~q ;
wire \D_logic_op_raw[1]~0_combout ;
wire \Equal154~2_combout ;
wire \Equal154~4_combout ;
wire \Equal154~5_combout ;
wire \D_ctrl_alu_force_xor~0_combout ;
wire \D_ctrl_alu_force_xor~1_combout ;
wire \D_ctrl_alu_force_xor~2_combout ;
wire \D_logic_op[1]~0_combout ;
wire \E_logic_op[1]~q ;
wire \D_logic_op_raw[0]~1_combout ;
wire \D_logic_op[0]~1_combout ;
wire \E_logic_op[0]~q ;
wire \E_logic_result[31]~9_combout ;
wire \E_alu_result~30_combout ;
wire \E_alu_result[31]~combout ;
wire \M_alu_result[31]~q ;
wire \E_op_rdctl~0_combout ;
wire \E_op_rdctl~combout ;
wire \M_ctrl_rdctl_inst~q ;
wire \M_ctrl_mem_nxt~0_combout ;
wire \M_ctrl_mem~q ;
wire \A_inst_result[31]~q ;
wire \D_ctrl_shift_rot~0_combout ;
wire \E_ctrl_shift_rot~q ;
wire \M_ctrl_shift_rot~q ;
wire \A_ctrl_shift_rot~q ;
wire \E_ld_bus~0_combout ;
wire \M_ctrl_ld_bypass~q ;
wire \A_ctrl_ld_bypass~q ;
wire \A_slow_inst_sel_nxt~0_combout ;
wire \A_slow_inst_sel~q ;
wire \E_ctrl_ld8_ld16~0_combout ;
wire \M_ctrl_ld8_ld16~q ;
wire \A_ld_align_byte2_byte3_fill~q ;
wire \A_wr_data_unfiltered[29]~32_combout ;
wire \A_mul_partial_prod[31]~q ;
wire \A_mul_partial_prod[30]~q ;
wire \A_mul_partial_prod[29]~q ;
wire \A_mul_partial_prod[28]~q ;
wire \A_mul_partial_prod[27]~q ;
wire \A_mul_partial_prod[26]~q ;
wire \A_mul_partial_prod[25]~q ;
wire \A_mul_partial_prod[24]~q ;
wire \A_mul_partial_prod[23]~q ;
wire \A_mul_partial_prod[22]~q ;
wire \A_mul_partial_prod[21]~q ;
wire \A_mul_partial_prod[20]~q ;
wire \A_mul_partial_prod[19]~q ;
wire \A_mul_partial_prod[18]~q ;
wire \A_mul_partial_prod[17]~q ;
wire \A_mul_partial_prod[16]~q ;
wire \A_mul_partial_prod[15]~q ;
wire \A_mul_partial_prod[14]~q ;
wire \A_mul_partial_prod[13]~q ;
wire \A_mul_partial_prod[12]~q ;
wire \A_mul_partial_prod[11]~q ;
wire \A_mul_partial_prod[10]~q ;
wire \A_mul_partial_prod[9]~q ;
wire \A_mul_partial_prod[8]~q ;
wire \A_mul_partial_prod[7]~q ;
wire \A_mul_partial_prod[6]~q ;
wire \A_mul_partial_prod[5]~q ;
wire \A_mul_partial_prod[4]~q ;
wire \A_mul_partial_prod[3]~q ;
wire \A_mul_partial_prod[2]~q ;
wire \A_mul_partial_prod[1]~q ;
wire \A_mul_partial_prod[0]~q ;
wire \Add19~53_sumout ;
wire \always120~0_combout ;
wire \A_mul_cnt_nxt[0]~2_combout ;
wire \A_mul_cnt[0]~q ;
wire \A_mul_cnt_nxt[1]~1_combout ;
wire \A_mul_cnt[1]~q ;
wire \A_mul_cnt_nxt[2]~0_combout ;
wire \A_mul_cnt[2]~q ;
wire \A_mul_stall_nxt~0_combout ;
wire \A_mul_stall~q ;
wire \A_mul_stall_d1~q ;
wire \A_mul_stall_d2~q ;
wire \A_mul_stall_d3~q ;
wire \A_mul_result[0]~q ;
wire \Add19~54 ;
wire \Add19~49_sumout ;
wire \A_mul_result[1]~q ;
wire \Add19~50 ;
wire \Add19~1_sumout ;
wire \A_mul_result[2]~q ;
wire \Add19~2 ;
wire \Add19~45_sumout ;
wire \A_mul_result[3]~q ;
wire \Add19~46 ;
wire \Add19~41_sumout ;
wire \A_mul_result[4]~q ;
wire \Add19~42 ;
wire \Add19~37_sumout ;
wire \A_mul_result[5]~q ;
wire \Add19~38 ;
wire \Add19~33_sumout ;
wire \A_mul_result[6]~q ;
wire \Add19~34 ;
wire \Add19~29_sumout ;
wire \A_mul_result[7]~q ;
wire \Add19~30 ;
wire \Add19~25_sumout ;
wire \A_mul_result[8]~q ;
wire \Add19~26 ;
wire \Add19~21_sumout ;
wire \A_mul_result[9]~q ;
wire \Add19~22 ;
wire \Add19~17_sumout ;
wire \A_mul_result[10]~q ;
wire \Add19~18 ;
wire \Add19~13_sumout ;
wire \A_mul_result[11]~q ;
wire \Add19~14 ;
wire \Add19~9_sumout ;
wire \A_mul_result[12]~q ;
wire \Add19~10 ;
wire \Add19~5_sumout ;
wire \A_mul_result[13]~q ;
wire \Add19~6 ;
wire \Add19~109_sumout ;
wire \A_mul_result[14]~q ;
wire \Add19~110 ;
wire \Add19~101_sumout ;
wire \A_mul_result[15]~q ;
wire \Add19~102 ;
wire \Add19~77_sumout ;
wire \A_mul_result[16]~q ;
wire \Add19~78 ;
wire \Add19~69_sumout ;
wire \A_mul_result[17]~q ;
wire \Add19~70 ;
wire \Add19~93_sumout ;
wire \A_mul_result[18]~q ;
wire \Add19~94 ;
wire \Add19~85_sumout ;
wire \A_mul_result[19]~q ;
wire \Add19~86 ;
wire \Add19~61_sumout ;
wire \A_mul_result[20]~q ;
wire \Add19~62 ;
wire \Add19~57_sumout ;
wire \A_mul_result[21]~q ;
wire \Add19~58 ;
wire \Add19~105_sumout ;
wire \A_mul_result[22]~q ;
wire \Add19~106 ;
wire \Add19~97_sumout ;
wire \A_mul_result[23]~q ;
wire \Add19~98 ;
wire \Add19~73_sumout ;
wire \A_mul_result[24]~q ;
wire \Add19~74 ;
wire \Add19~65_sumout ;
wire \A_mul_result[25]~q ;
wire \Add19~66 ;
wire \Add19~89_sumout ;
wire \A_mul_result[26]~q ;
wire \Add19~90 ;
wire \Add19~81_sumout ;
wire \A_mul_result[27]~q ;
wire \Add19~82 ;
wire \Add19~125_sumout ;
wire \A_mul_result[28]~q ;
wire \Add19~126 ;
wire \Add19~113_sumout ;
wire \A_mul_result[29]~q ;
wire \Add19~114 ;
wire \Add19~117_sumout ;
wire \A_mul_result[30]~q ;
wire \Add19~118 ;
wire \Add19~121_sumout ;
wire \A_mul_result[31]~q ;
wire \D_iw[6]~q ;
wire \E_compare_op[0]~q ;
wire \D_src2_reg[0]~28_combout ;
wire \E_alu_result~20_combout ;
wire \E_alu_result[27]~combout ;
wire \M_alu_result[27]~q ;
wire \A_inst_result[27]~q ;
wire \E_ctrl_ld_signed~0_combout ;
wire \M_ctrl_ld_signed~q ;
wire \A_ctrl_ld_signed~q ;
wire \D_ctrl_shift_right_arith~0_combout ;
wire \D_ctrl_shift_right_arith~1_combout ;
wire \E_ctrl_shift_right_arith~q ;
wire \E_rot_fill_bit~0_combout ;
wire \M_rot_fill_bit~q ;
wire \D_iw[8]~q ;
wire \d_readdata_d1[2]~q ;
wire \d_readdata_d1[10]~q ;
wire \d_readdata_d1[18]~q ;
wire \d_readdata_d1[26]~q ;
wire \M_alu_result[0]~q ;
wire \Equal184~0_combout ;
wire \M_ctrl_ld8~q ;
wire \M_ld_align_sh8~0_combout ;
wire \A_ld_align_sh8~q ;
wire \D_iw[7]~q ;
wire \D_src2_reg[5]~3_combout ;
wire \D_src2_reg[5]~4_combout ;
wire \d_readdata_d1[1]~q ;
wire \d_readdata_d1[9]~q ;
wire \d_readdata_d1[17]~q ;
wire \d_readdata_d1[25]~q ;
wire \A_slow_ld_byte0_data_aligned_nxt[1]~6_combout ;
wire \d_readdatavalid_d1~q ;
wire \D_iw[10]~q ;
wire \d_readdata_d1[4]~q ;
wire \d_readdata_d1[12]~q ;
wire \d_readdata_d1[20]~q ;
wire \d_readdata_d1[28]~q ;
wire \A_slow_ld_byte0_data_aligned_nxt[4]~4_combout ;
wire \A_slow_inst_result[4]~q ;
wire \A_inst_result[4]~q ;
wire \D_src2_reg[13]~8_combout ;
wire \D_iw[9]~q ;
wire \d_readdata_d1[3]~q ;
wire \d_readdata_d1[11]~q ;
wire \d_readdata_d1[19]~q ;
wire \d_readdata_d1[27]~q ;
wire \A_slow_ld_byte0_data_aligned_nxt[3]~5_combout ;
wire \A_slow_inst_result[3]~q ;
wire \A_inst_result[3]~q ;
wire \E_ctrl_shift_rot_right~q ;
wire \D_ctrl_shift_rot_left~0_combout ;
wire \E_ctrl_shift_rot_left~q ;
wire \E_rot_sel_fill1~0_combout ;
wire \M_rot_sel_fill1~q ;
wire \d_readdata_d1[7]~q ;
wire \d_readdata_d1[15]~q ;
wire \d_readdata_d1[23]~q ;
wire \d_readdata_d1[31]~q ;
wire \A_slow_ld_byte0_data_aligned_nxt[7]~1_combout ;
wire \A_slow_inst_result[7]~q ;
wire \D_src2_reg[7]~14_combout ;
wire \D_src2_reg[7]~15_combout ;
wire \F_ctrl_hi_imm16~0_combout ;
wire \D_ctrl_hi_imm16~q ;
wire \E_src2[14]~0_combout ;
wire \E_src2[7]~q ;
wire \d_readdata_d1[6]~q ;
wire \d_readdata_d1[14]~q ;
wire \d_readdata_d1[22]~q ;
wire \d_readdata_d1[30]~q ;
wire \A_slow_ld_byte0_data_aligned_nxt[6]~2_combout ;
wire \A_slow_inst_result[6]~q ;
wire \A_inst_result[6]~q ;
wire \E_rot_mask[6]~7_combout ;
wire \M_rot_mask[6]~q ;
wire \E_rot_mask[2]~0_combout ;
wire \M_rot_mask[2]~q ;
wire \d_readdata_d1[5]~q ;
wire \d_readdata_d1[13]~q ;
wire \d_readdata_d1[21]~q ;
wire \d_readdata_d1[29]~q ;
wire \A_slow_ld_byte0_data_aligned_nxt[5]~3_combout ;
wire \A_slow_inst_result[5]~q ;
wire \D_src2_reg[5]~18_combout ;
wire \D_src2_reg[5]~19_combout ;
wire \E_src2[5]~q ;
wire \E_regnum_a_cmp_F~0_combout ;
wire \E_regnum_a_cmp_F~1_combout ;
wire \E_regnum_a_cmp_F~combout ;
wire \D_regnum_a_cmp_F~0_combout ;
wire \D_regnum_a_cmp_F~combout ;
wire \E_regnum_a_cmp_D~q ;
wire \M_regnum_a_cmp_D~q ;
wire \A_regnum_a_cmp_F~0_combout ;
wire \A_regnum_a_cmp_F~1_combout ;
wire \A_regnum_a_cmp_F~combout ;
wire \M_regnum_a_cmp_F~0_combout ;
wire \M_regnum_a_cmp_F~1_combout ;
wire \M_regnum_a_cmp_F~combout ;
wire \A_regnum_a_cmp_D~q ;
wire \W_regnum_a_cmp_D~q ;
wire \E_src1[7]~0_combout ;
wire \E_src1[7]~1_combout ;
wire \D_src1_reg[4]~10_combout ;
wire \D_iw[28]~q ;
wire \D_iw[29]~q ;
wire \D_iw[31]~q ;
wire \D_iw[30]~q ;
wire \D_iw[27]~q ;
wire \Equal296~0_combout ;
wire \D_src1_hazard_E~combout ;
wire \E_src1[4]~q ;
wire \D_src1_reg[1]~30_combout ;
wire \E_src1[1]~q ;
wire \d_readdata_d1[0]~q ;
wire \d_readdata_d1[8]~q ;
wire \d_readdata_d1[16]~q ;
wire \d_readdata_d1[24]~q ;
wire \A_slow_ld_byte0_data_aligned_nxt[0]~7_combout ;
wire \A_slow_inst_result[0]~q ;
wire \M_inst_result~0_combout ;
wire \D_ctrl_crst~0_combout ;
wire \E_ctrl_crst~q ;
wire \M_ctrl_crst~q ;
wire \D_ctrl_break~0_combout ;
wire \E_ctrl_break~q ;
wire \M_ctrl_break~q ;
wire \D_ctrl_exception~0_combout ;
wire \E_ctrl_exception~q ;
wire \M_ctrl_exception~q ;
wire \M_iw[14]~q ;
wire \M_iw[11]~q ;
wire \M_iw[5]~q ;
wire \M_iw[0]~q ;
wire \M_iw[16]~q ;
wire \M_iw[15]~q ;
wire \M_iw[13]~q ;
wire \M_iw[12]~q ;
wire \M_op_eret~0_combout ;
wire \M_iw[4]~q ;
wire \M_iw[3]~q ;
wire \M_iw[2]~q ;
wire \M_iw[1]~q ;
wire \M_op_eret~1_combout ;
wire \M_op_eret~2_combout ;
wire \E_iw[6]~q ;
wire \M_iw[6]~q ;
wire \E_iw[7]~q ;
wire \M_iw[7]~q ;
wire \E_iw[8]~q ;
wire \M_iw[8]~q ;
wire \E_op_wrctl~combout ;
wire \M_ctrl_wrctl_inst~q ;
wire \M_wrctl_bstatus~combout ;
wire \A_bstatus_reg_pie_inst_nxt~0_combout ;
wire \A_bstatus_reg_pie~q ;
wire \A_status_reg_pie_inst_nxt~0_combout ;
wire \A_status_reg_pie_inst_nxt~1_combout ;
wire \A_status_reg_pie_inst_nxt~2_combout ;
wire \A_status_reg_pie~q ;
wire \M_wrctl_estatus~combout ;
wire \A_estatus_reg_pie_inst_nxt~0_combout ;
wire \A_estatus_reg_pie~q ;
wire \D_control_reg_rddata_muxed[0]~0_combout ;
wire \E_control_reg_rddata[0]~q ;
wire \M_control_reg_rddata[0]~q ;
wire \A_inst_result[0]~q ;
wire \E_rot_mask[0]~5_combout ;
wire \M_rot_mask[0]~q ;
wire \Add7~0_combout ;
wire \E_rot_step1[4]~19_combout ;
wire \D_src1_reg[8]~6_combout ;
wire \E_src1[8]~q ;
wire \E_rot_step1[8]~16_combout ;
wire \Add7~1_combout ;
wire \M_rot_prestep2[8]~q ;
wire \D_src1_reg[17]~16_combout ;
wire \E_src1[17]~q ;
wire \E_alu_result~17_combout ;
wire \D_src1_reg[16]~17_combout ;
wire \E_src1[16]~q ;
wire \E_alu_result~19_combout ;
wire \E_rot_mask[7]~6_combout ;
wire \M_rot_mask[7]~q ;
wire \D_src1_reg[11]~3_combout ;
wire \E_src1[11]~q ;
wire \E_rot_mask[1]~4_combout ;
wire \M_rot_mask[1]~q ;
wire \E_rot_step1[5]~11_combout ;
wire \E_rot_step1[9]~8_combout ;
wire \M_rot_prestep2[9]~q ;
wire \Add17~134 ;
wire \Add17~129_sumout ;
wire \D_src2_reg[29]~57_combout ;
wire \D_src2_reg[29]~58_combout ;
wire \F_ctrl_unsigned_lo_imm16~1_combout ;
wire \F_ctrl_unsigned_lo_imm16~0_combout ;
wire \D_ctrl_unsigned_lo_imm16~q ;
wire \D_src2[29]~2_combout ;
wire \D_src2[29]~3_combout ;
wire \E_src2[19]~1_combout ;
wire \E_src2[29]~q ;
wire \E_logic_result[29]~7_combout ;
wire \E_alu_result~28_combout ;
wire \E_alu_result[29]~combout ;
wire \M_alu_result[29]~q ;
wire \A_inst_result[29]~q ;
wire \E_rot_mask[5]~1_combout ;
wire \M_rot_mask[5]~q ;
wire \D_ctrl_rot~0_combout ;
wire \E_ctrl_rot~q ;
wire \E_rot_pass3~0_combout ;
wire \M_rot_pass3~q ;
wire \E_rot_sel_fill3~0_combout ;
wire \M_rot_sel_fill3~q ;
wire \E_rot_step1[25]~12_combout ;
wire \M_rot_prestep2[29]~q ;
wire \D_src1_reg[14]~27_combout ;
wire \E_src1[14]~q ;
wire \E_rot_step1[17]~14_combout ;
wire \E_rot_step1[21]~15_combout ;
wire \M_rot_prestep2[21]~q ;
wire \E_logic_result[30]~8_combout ;
wire \E_alu_result~29_combout ;
wire \D_src2_reg[30]~59_combout ;
wire \D_src2_reg[30]~60_combout ;
wire \D_src2[30]~4_combout ;
wire \D_src2[30]~5_combout ;
wire \E_src2[30]~q ;
wire \Add17~130 ;
wire \Add17~65_sumout ;
wire \E_alu_result[30]~combout ;
wire \M_alu_result[30]~q ;
wire \A_inst_result[30]~q ;
wire \E_rot_step1[26]~3_combout ;
wire \E_rot_step1[30]~0_combout ;
wire \M_rot_prestep2[30]~q ;
wire \E_rot_step1[18]~5_combout ;
wire \E_rot_step1[22]~2_combout ;
wire \M_rot_prestep2[22]~q ;
wire \E_rot_step1[2]~1_combout ;
wire \M_rot_prestep2[6]~q ;
wire \Add7~2_combout ;
wire \M_rot_rn[3]~q ;
wire \Add7~3_combout ;
wire \M_rot_rn[4]~q ;
wire \M_rot[6]~29_combout ;
wire \A_shift_rot_result~29_combout ;
wire \A_shift_rot_result[30]~q ;
wire \A_mem_baddr[1]~q ;
wire \A_mem_baddr[0]~q ;
wire \Equal187~0_combout ;
wire \M_ctrl_ld16~q ;
wire \A_ctrl_ld16~q ;
wire \A_slow_ld_data_sign_bit~0_combout ;
wire \A_slow_ld_data_fill_bit~0_combout ;
wire \A_slow_inst_result[30]~q ;
wire \A_wr_data_unfiltered[30]~61_combout ;
wire \A_wr_data_unfiltered[30]~62_combout ;
wire \W_wr_data[30]~q ;
wire \D_src1_reg[30]~14_combout ;
wire \E_src1[30]~q ;
wire \E_rot_step1[1]~10_combout ;
wire \M_rot_prestep2[5]~q ;
wire \M_rot[5]~1_combout ;
wire \A_shift_rot_result~1_combout ;
wire \A_shift_rot_result[13]~q ;
wire \D_src2_reg[13]~7_combout ;
wire \D_src2_reg[13]~92_combout ;
wire \E_logic_result[13]~0_combout ;
wire \E_ctrl_jmp_indirect_nxt~0_combout ;
wire \E_valid_jmp_indirect~0_combout ;
wire \E_valid_jmp_indirect~q ;
wire \D_pc[11]~q ;
wire \D_src1_reg[12]~2_combout ;
wire \E_src1[12]~q ;
wire \D_pc[10]~q ;
wire \Add3~1_sumout ;
wire \Add0~1_sumout ;
wire \D_br_taken_waddr_partial[0]~q ;
wire \D_pc_plus_one[0]~q ;
wire \E_ctrl_br_cond_nxt~0_combout ;
wire \D_br_pred_not_taken~combout ;
wire \E_extra_pc[0]~q ;
wire \E_ctrl_jmp_indirect~q ;
wire \M_pipe_flush_waddr[0]~0_combout ;
wire \M_pipe_flush_waddr_nxt[0]~0_combout ;
wire \D_pc[0]~q ;
wire \E_pc[0]~q ;
wire \M_pipe_flush_waddr[0]~1_combout ;
wire \M_pipe_flush_waddr[0]~q ;
wire \D_kill~q ;
wire \F_ctrl_br~0_combout ;
wire \D_ctrl_br~q ;
wire \F_ctrl_br_uncond~0_combout ;
wire \D_ctrl_br_uncond~q ;
wire \F_ic_data_rd_addr_nxt[2]~1_combout ;
wire \F_ic_data_rd_addr_nxt[0]~2_combout ;
wire \F_ic_data_rd_addr_nxt[0]~3_combout ;
wire \F_pc[0]~q ;
wire \Add3~2 ;
wire \Add3~45_sumout ;
wire \Add0~2 ;
wire \Add0~41_sumout ;
wire \D_br_taken_waddr_partial[1]~q ;
wire \D_pc_plus_one[1]~q ;
wire \E_extra_pc[1]~q ;
wire \M_pipe_flush_waddr_nxt[1]~1_combout ;
wire \D_pc[1]~q ;
wire \E_pc[1]~q ;
wire \M_pipe_flush_waddr[1]~q ;
wire \F_ic_data_rd_addr_nxt[1]~4_combout ;
wire \F_ic_data_rd_addr_nxt[1]~5_combout ;
wire \F_pc[1]~q ;
wire \Add3~46 ;
wire \Add3~41_sumout ;
wire \Add0~42 ;
wire \Add0~37_sumout ;
wire \D_br_taken_waddr_partial[2]~q ;
wire \D_pc_plus_one[2]~q ;
wire \E_extra_pc[2]~q ;
wire \M_pipe_flush_waddr_nxt[2]~2_combout ;
wire \D_pc[2]~q ;
wire \E_pc[2]~q ;
wire \M_pipe_flush_waddr[2]~q ;
wire \F_ic_data_rd_addr_nxt[2]~6_combout ;
wire \F_ic_data_rd_addr_nxt[2]~7_combout ;
wire \F_pc[2]~q ;
wire \Add3~42 ;
wire \Add3~37_sumout ;
wire \Add0~38 ;
wire \Add0~33_sumout ;
wire \D_br_taken_waddr_partial[3]~q ;
wire \D_pc_plus_one[3]~q ;
wire \E_extra_pc[3]~q ;
wire \M_pipe_flush_waddr_nxt[3]~3_combout ;
wire \D_pc[3]~q ;
wire \E_pc[3]~q ;
wire \M_pipe_flush_waddr[3]~q ;
wire \F_ic_tag_rd_addr_nxt[0]~0_combout ;
wire \F_ic_tag_rd_addr_nxt[0]~1_combout ;
wire \F_pc[3]~q ;
wire \Add3~38 ;
wire \Add3~33_sumout ;
wire \Add0~34 ;
wire \Add0~29_sumout ;
wire \D_br_taken_waddr_partial[4]~q ;
wire \D_pc_plus_one[4]~q ;
wire \E_extra_pc[4]~q ;
wire \M_pipe_flush_waddr_nxt[4]~4_combout ;
wire \D_pc[4]~q ;
wire \E_pc[4]~q ;
wire \M_pipe_flush_waddr[4]~q ;
wire \F_ic_tag_rd_addr_nxt[1]~2_combout ;
wire \F_ic_tag_rd_addr_nxt[1]~3_combout ;
wire \F_pc[4]~q ;
wire \Add3~34 ;
wire \Add3~29_sumout ;
wire \Add0~30 ;
wire \Add0~25_sumout ;
wire \D_br_taken_waddr_partial[5]~q ;
wire \D_pc_plus_one[5]~q ;
wire \E_extra_pc[5]~q ;
wire \M_pipe_flush_waddr_nxt[5]~5_combout ;
wire \D_pc[5]~q ;
wire \E_pc[5]~q ;
wire \M_pipe_flush_waddr[5]~q ;
wire \F_ic_tag_rd_addr_nxt[2]~4_combout ;
wire \F_ic_tag_rd_addr_nxt[2]~5_combout ;
wire \F_pc[5]~q ;
wire \Add3~30 ;
wire \Add3~25_sumout ;
wire \Add0~26 ;
wire \Add0~21_sumout ;
wire \D_br_taken_waddr_partial[6]~q ;
wire \D_pc_plus_one[6]~q ;
wire \E_extra_pc[6]~q ;
wire \M_pipe_flush_waddr_nxt[6]~6_combout ;
wire \D_pc[6]~q ;
wire \E_pc[6]~q ;
wire \M_pipe_flush_waddr[6]~q ;
wire \F_ic_tag_rd_addr_nxt[3]~6_combout ;
wire \F_ic_tag_rd_addr_nxt[3]~7_combout ;
wire \F_pc[6]~q ;
wire \Add3~26 ;
wire \Add3~21_sumout ;
wire \Add0~22 ;
wire \Add0~17_sumout ;
wire \D_br_taken_waddr_partial[7]~q ;
wire \D_pc_plus_one[7]~q ;
wire \E_extra_pc[7]~q ;
wire \M_pipe_flush_waddr_nxt[7]~7_combout ;
wire \D_pc[7]~q ;
wire \E_pc[7]~q ;
wire \M_pipe_flush_waddr[7]~q ;
wire \F_ic_tag_rd_addr_nxt[4]~8_combout ;
wire \F_ic_tag_rd_addr_nxt[4]~9_combout ;
wire \F_pc[7]~q ;
wire \Add3~22 ;
wire \Add3~17_sumout ;
wire \Add0~18 ;
wire \Add0~13_sumout ;
wire \D_br_taken_waddr_partial[8]~q ;
wire \D_pc_plus_one[8]~q ;
wire \E_extra_pc[8]~q ;
wire \M_pipe_flush_waddr_nxt[8]~8_combout ;
wire \D_pc[8]~q ;
wire \E_pc[8]~q ;
wire \M_pipe_flush_waddr[8]~q ;
wire \F_ic_tag_rd_addr_nxt[5]~10_combout ;
wire \F_ic_tag_rd_addr_nxt[5]~11_combout ;
wire \F_pc[8]~q ;
wire \Add3~18 ;
wire \Add3~13_sumout ;
wire \Add0~14 ;
wire \Add0~9_sumout ;
wire \D_br_taken_waddr_partial[9]~q ;
wire \D_pc_plus_one[9]~q ;
wire \E_extra_pc[9]~q ;
wire \M_pipe_flush_waddr_nxt[9]~9_combout ;
wire \D_pc[9]~q ;
wire \E_pc[9]~q ;
wire \M_pipe_flush_waddr[9]~q ;
wire \F_ic_tag_rd_addr_nxt[6]~12_combout ;
wire \F_ic_tag_rd_addr_nxt[6]~13_combout ;
wire \F_pc[9]~q ;
wire \Add3~14 ;
wire \Add3~9_sumout ;
wire \D_pc_plus_one[10]~q ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \D_br_taken_waddr_partial[10]~q ;
wire \Add1~1_combout ;
wire \F_pc_nxt~0_combout ;
wire \F_pc_nxt~1_combout ;
wire \E_pc[10]~q ;
wire \E_extra_pc[10]~q ;
wire \M_pipe_flush_waddr_nxt[10]~10_combout ;
wire \M_pipe_flush_waddr_nxt[10]~11_combout ;
wire \M_pipe_flush_waddr[10]~q ;
wire \M_pipe_flush_waddr[10]~_wirecell_combout ;
wire \F_pc[10]~q ;
wire \F_ic_valid~4_combout ;
wire \F_ic_valid~0_combout ;
wire \F_ic_hit~0_combout ;
wire \D_iw_valid~q ;
wire \D_br_pred_taken~0_combout ;
wire \F_kill~2_combout ;
wire \F_kill~0_combout ;
wire \F_kill~1_combout ;
wire \F_issue~combout ;
wire \D_issue~q ;
wire \F_ic_data_rd_addr_nxt[2]~0_combout ;
wire \F_pc_nxt~2_combout ;
wire \F_pc_nxt~3_combout ;
wire \M_pipe_flush_waddr_nxt[11]~12_combout ;
wire \E_pc[11]~q ;
wire \M_pipe_flush_waddr[11]~q ;
wire \F_pc[11]~q ;
wire \Add3~10 ;
wire \Add3~5_sumout ;
wire \D_pc_plus_one[11]~q ;
wire \Add1~0_combout ;
wire \E_extra_pc[11]~q ;
wire \E_alu_result[13]~2_combout ;
wire \D_src2_reg[13]~128_combout ;
wire \E_src2[13]~q ;
wire \Add17~10 ;
wire \Add17~2 ;
wire \Add17~5_sumout ;
wire \E_logic_result[9]~4_combout ;
wire \E_alu_result[9]~6_combout ;
wire \E_alu_result[9]~combout ;
wire \M_alu_result[9]~q ;
wire \A_inst_result[9]~q ;
wire \A_ld_align_byte1_fill~q ;
wire \A_slow_ld_byte1_data_aligned_nxt[1]~4_combout ;
wire \A_slow_inst_result[9]~q ;
wire \A_data_ram_ld_align_fill_bit~combout ;
wire \A_wr_data_unfiltered[11]~4_combout ;
wire \A_wr_data_unfiltered[11]~5_combout ;
wire \A_wr_data_unfiltered[9]~14_combout ;
wire \D_src2_reg[9]~12_combout ;
wire \D_src2_reg[9]~96_combout ;
wire \D_src2_reg[9]~112_combout ;
wire \E_src2[9]~q ;
wire \Add17~6 ;
wire \Add17~13_sumout ;
wire \E_logic_result[10]~3_combout ;
wire \E_alu_result[10]~5_combout ;
wire \E_alu_result[10]~combout ;
wire \M_alu_result[10]~q ;
wire \A_inst_result[10]~q ;
wire \A_slow_ld_byte1_data_aligned_nxt[2]~3_combout ;
wire \A_slow_inst_result[10]~q ;
wire \A_wr_data_unfiltered[10]~12_combout ;
wire \D_src2_reg[10]~11_combout ;
wire \D_src2_reg[10]~95_combout ;
wire \D_src2_reg[10]~116_combout ;
wire \E_src2[10]~q ;
wire \Add17~14 ;
wire \Add17~50 ;
wire \Add17~46 ;
wire \Add17~41_sumout ;
wire \E_alu_result[13]~combout ;
wire \M_alu_result[13]~q ;
wire \A_inst_result[13]~q ;
wire \A_slow_ld_byte1_data_aligned_nxt[5]~0_combout ;
wire \A_slow_inst_result[13]~q ;
wire \A_wr_data_unfiltered[13]~6_combout ;
wire \A_wr_data_unfiltered[13]~7_combout ;
wire \W_wr_data[13]~q ;
wire \D_src1_reg[13]~1_combout ;
wire \E_src1[13]~q ;
wire \E_rot_step1[13]~9_combout ;
wire \M_rot_prestep2[13]~q ;
wire \M_rot[5]~28_combout ;
wire \A_shift_rot_result~28_combout ;
wire \A_shift_rot_result[29]~q ;
wire \A_slow_inst_result[29]~q ;
wire \A_wr_data_unfiltered[29]~59_combout ;
wire \A_wr_data_unfiltered[29]~60_combout ;
wire \W_wr_data[29]~q ;
wire \D_src1_reg[29]~13_combout ;
wire \E_src1[29]~q ;
wire \E_rot_step1[29]~13_combout ;
wire \M_rot_prestep2[1]~q ;
wire \M_rot_prestep2[25]~q ;
wire \M_rot_prestep2[17]~q ;
wire \M_rot[1]~5_combout ;
wire \A_shift_rot_result~5_combout ;
wire \A_shift_rot_result[9]~q ;
wire \A_wr_data_unfiltered[9]~15_combout ;
wire \W_wr_data[9]~q ;
wire \D_src1_reg[9]~5_combout ;
wire \E_src1[9]~q ;
wire \E_rot_step1[11]~25_combout ;
wire \E_rot_step1[15]~30_combout ;
wire \M_rot_prestep2[15]~q ;
wire \E_rot_step1[3]~27_combout ;
wire \M_rot_prestep2[7]~q ;
wire \E_rot_step1[27]~29_combout ;
wire \E_rot_step1[31]~26_combout ;
wire \M_rot_prestep2[31]~q ;
wire \E_rot_step1[19]~31_combout ;
wire \E_rot_step1[23]~28_combout ;
wire \M_rot_prestep2[23]~q ;
wire \M_rot[7]~25_combout ;
wire \A_shift_rot_result~25_combout ;
wire \A_shift_rot_result[15]~q ;
wire \A_inst_result[15]~q ;
wire \A_slow_ld_byte1_data_aligned_nxt[7]~6_combout ;
wire \A_slow_inst_result[15]~q ;
wire \A_wr_data_unfiltered[15]~55_combout ;
wire \A_wr_data_unfiltered[15]~67_combout ;
wire \W_wr_data[15]~q ;
wire \D_src1_reg[15]~23_combout ;
wire \E_src1[15]~q ;
wire \E_logic_result[15]~11_combout ;
wire \E_alu_result~25_combout ;
wire \Add17~42 ;
wire \Add17~126 ;
wire \Add17~117_sumout ;
wire \E_alu_result[15]~combout ;
wire \M_alu_result[15]~q ;
wire \D_src2_reg[15]~51_combout ;
wire \D_src2_reg[15]~98_combout ;
wire \D_src2_reg[15]~104_combout ;
wire \E_src2[15]~q ;
wire \Add17~118 ;
wire \Add17~93_sumout ;
wire \E_alu_result[16]~combout ;
wire \M_alu_result[16]~q ;
wire \A_inst_result[16]~q ;
wire \E_rot_pass2~0_combout ;
wire \M_rot_pass2~q ;
wire \E_rot_sel_fill2~0_combout ;
wire \M_rot_sel_fill2~q ;
wire \E_rot_step1[12]~17_combout ;
wire \E_rot_step1[16]~22_combout ;
wire \M_rot_prestep2[16]~q ;
wire \E_rot_step1[20]~23_combout ;
wire \E_rot_step1[24]~20_combout ;
wire \M_rot_prestep2[24]~q ;
wire \M_rot[0]~19_combout ;
wire \A_shift_rot_result~19_combout ;
wire \A_shift_rot_result[16]~q ;
wire \A_slow_inst_result[16]~q ;
wire \A_wr_data_unfiltered[16]~43_combout ;
wire \A_wr_data_unfiltered[16]~44_combout ;
wire \W_wr_data[16]~q ;
wire \D_src2_reg[16]~39_combout ;
wire \D_src2[16]~32_combout ;
wire \D_src2[16]~33_combout ;
wire \D_src2[16]~9_combout ;
wire \E_src2[16]~q ;
wire \Add17~94 ;
wire \Add17~85_sumout ;
wire \E_alu_result[17]~combout ;
wire \M_alu_result[17]~q ;
wire \A_inst_result[17]~q ;
wire \M_rot[1]~17_combout ;
wire \A_shift_rot_result~17_combout ;
wire \A_shift_rot_result[17]~q ;
wire \A_slow_inst_result[17]~q ;
wire \A_wr_data_unfiltered[17]~39_combout ;
wire \A_wr_data_unfiltered[17]~40_combout ;
wire \W_wr_data[17]~q ;
wire \D_src2_reg[17]~35_combout ;
wire \D_src2[17]~30_combout ;
wire \D_src2[17]~31_combout ;
wire \D_src2[17]~8_combout ;
wire \E_src2[17]~q ;
wire \Add17~86 ;
wire \Add17~109_sumout ;
wire \E_alu_result[18]~combout ;
wire \M_alu_result[18]~q ;
wire \A_inst_result[18]~q ;
wire \E_rot_step1[14]~4_combout ;
wire \M_rot_prestep2[18]~q ;
wire \M_rot_prestep2[2]~q ;
wire \M_rot_prestep2[26]~q ;
wire \M_rot[2]~23_combout ;
wire \A_shift_rot_result~23_combout ;
wire \A_shift_rot_result[18]~q ;
wire \A_slow_inst_result[18]~q ;
wire \A_wr_data_unfiltered[18]~51_combout ;
wire \A_wr_data_unfiltered[18]~52_combout ;
wire \W_wr_data[18]~q ;
wire \D_src1_reg[18]~19_combout ;
wire \E_src1[18]~q ;
wire \E_alu_result~23_combout ;
wire \D_src2_reg[18]~65_combout ;
wire \D_src2_reg[18]~47_combout ;
wire \D_src2[18]~12_combout ;
wire \D_src2[18]~13_combout ;
wire \E_src2[18]~q ;
wire \Add17~110 ;
wire \Add17~101_sumout ;
wire \E_alu_result[19]~combout ;
wire \M_alu_result[19]~q ;
wire \A_inst_result[19]~q ;
wire \M_rot_prestep2[19]~q ;
wire \M_rot_prestep2[3]~q ;
wire \M_rot_prestep2[27]~q ;
wire \M_rot[3]~21_combout ;
wire \A_shift_rot_result~21_combout ;
wire \A_shift_rot_result[19]~q ;
wire \A_slow_inst_result[19]~q ;
wire \A_wr_data_unfiltered[19]~47_combout ;
wire \A_wr_data_unfiltered[19]~48_combout ;
wire \W_wr_data[19]~q ;
wire \D_src1_reg[19]~21_combout ;
wire \E_src1[19]~q ;
wire \E_alu_result~21_combout ;
wire \D_src2_reg[19]~67_combout ;
wire \D_src2_reg[19]~43_combout ;
wire \D_src2[19]~16_combout ;
wire \D_src2[19]~17_combout ;
wire \E_src2[19]~q ;
wire \Add17~102 ;
wire \Add17~77_sumout ;
wire \E_alu_result[20]~combout ;
wire \M_alu_result[20]~q ;
wire \A_inst_result[20]~q ;
wire \E_rot_mask[4]~2_combout ;
wire \M_rot_mask[4]~q ;
wire \M_rot_prestep2[20]~q ;
wire \M_rot_prestep2[12]~q ;
wire \E_rot_step1[0]~18_combout ;
wire \M_rot_prestep2[4]~q ;
wire \M_rot_prestep2[28]~q ;
wire \M_rot[4]~15_combout ;
wire \A_shift_rot_result~15_combout ;
wire \A_shift_rot_result[20]~q ;
wire \A_slow_inst_result[20]~q ;
wire \A_wr_data_unfiltered[20]~35_combout ;
wire \A_wr_data_unfiltered[20]~36_combout ;
wire \W_wr_data[20]~q ;
wire \D_src1_reg[20]~25_combout ;
wire \E_src1[20]~q ;
wire \E_alu_result~15_combout ;
wire \D_src2_reg[20]~70_combout ;
wire \D_src2_reg[20]~31_combout ;
wire \D_src2[20]~22_combout ;
wire \D_src2[20]~23_combout ;
wire \E_src2[20]~q ;
wire \Add17~78 ;
wire \Add17~73_sumout ;
wire \E_alu_result[21]~combout ;
wire \M_alu_result[21]~q ;
wire \A_inst_result[21]~q ;
wire \M_rot[5]~14_combout ;
wire \A_shift_rot_result~14_combout ;
wire \A_shift_rot_result[21]~q ;
wire \A_slow_inst_result[21]~q ;
wire \A_wr_data_unfiltered[21]~33_combout ;
wire \A_wr_data_unfiltered[21]~34_combout ;
wire \W_wr_data[21]~q ;
wire \D_src1_reg[21]~22_combout ;
wire \E_src1[21]~q ;
wire \E_logic_result[21]~10_combout ;
wire \E_alu_result~14_combout ;
wire \D_src2_reg[21]~68_combout ;
wire \D_src2_reg[21]~29_combout ;
wire \D_src2[21]~18_combout ;
wire \D_src2[21]~19_combout ;
wire \E_src2[21]~q ;
wire \Add17~74 ;
wire \Add17~121_sumout ;
wire \E_alu_result[22]~combout ;
wire \M_alu_result[22]~q ;
wire \A_inst_result[22]~q ;
wire \M_rot[6]~26_combout ;
wire \A_shift_rot_result~26_combout ;
wire \A_shift_rot_result[22]~q ;
wire \A_slow_inst_result[22]~q ;
wire \A_wr_data_unfiltered[22]~56_combout ;
wire \A_wr_data_unfiltered[22]~57_combout ;
wire \W_wr_data[22]~q ;
wire \D_src1_reg[22]~26_combout ;
wire \E_src1[22]~q ;
wire \E_alu_result~26_combout ;
wire \D_src2_reg[22]~71_combout ;
wire \D_src2_reg[22]~52_combout ;
wire \D_src2[22]~24_combout ;
wire \D_src2[22]~25_combout ;
wire \E_src2[22]~q ;
wire \Add17~122 ;
wire \Add17~113_sumout ;
wire \E_alu_result[23]~combout ;
wire \M_alu_result[23]~q ;
wire \A_inst_result[23]~q ;
wire \M_rot[7]~24_combout ;
wire \A_shift_rot_result~24_combout ;
wire \A_shift_rot_result[23]~q ;
wire \A_slow_inst_result[23]~q ;
wire \A_wr_data_unfiltered[23]~53_combout ;
wire \A_wr_data_unfiltered[23]~54_combout ;
wire \W_wr_data[23]~q ;
wire \D_src1_reg[23]~29_combout ;
wire \E_src1[23]~q ;
wire \E_alu_result~24_combout ;
wire \D_src2_reg[23]~73_combout ;
wire \D_src2_reg[23]~49_combout ;
wire \D_src2[23]~28_combout ;
wire \D_src2[23]~29_combout ;
wire \E_src2[23]~q ;
wire \Add17~114 ;
wire \Add17~89_sumout ;
wire \E_alu_result[24]~combout ;
wire \M_alu_result[24]~q ;
wire \A_inst_result[24]~q ;
wire \M_rot[0]~18_combout ;
wire \A_shift_rot_result~18_combout ;
wire \A_shift_rot_result[24]~q ;
wire \A_slow_inst_result[24]~q ;
wire \A_wr_data_unfiltered[24]~41_combout ;
wire \A_wr_data_unfiltered[24]~42_combout ;
wire \W_wr_data[24]~q ;
wire \D_src1_reg[24]~28_combout ;
wire \E_src1[24]~q ;
wire \E_alu_result~18_combout ;
wire \D_src2_reg[24]~72_combout ;
wire \D_src2_reg[24]~37_combout ;
wire \D_src2[24]~26_combout ;
wire \D_src2[24]~27_combout ;
wire \E_src2[24]~q ;
wire \Add17~90 ;
wire \Add17~81_sumout ;
wire \E_alu_result[25]~combout ;
wire \M_alu_result[25]~q ;
wire \A_inst_result[25]~q ;
wire \M_rot[1]~16_combout ;
wire \A_shift_rot_result~16_combout ;
wire \A_shift_rot_result[25]~q ;
wire \A_slow_inst_result[25]~q ;
wire \A_wr_data_unfiltered[25]~37_combout ;
wire \A_wr_data_unfiltered[25]~38_combout ;
wire \W_wr_data[25]~q ;
wire \D_src1_reg[25]~24_combout ;
wire \E_src1[25]~q ;
wire \E_alu_result~16_combout ;
wire \D_src2_reg[25]~69_combout ;
wire \D_src2_reg[25]~33_combout ;
wire \D_src2[25]~20_combout ;
wire \D_src2[25]~21_combout ;
wire \E_src2[25]~q ;
wire \Add17~82 ;
wire \Add17~105_sumout ;
wire \E_alu_result[26]~combout ;
wire \M_alu_result[26]~q ;
wire \A_inst_result[26]~q ;
wire \M_rot[2]~22_combout ;
wire \A_shift_rot_result~22_combout ;
wire \A_shift_rot_result[26]~q ;
wire \A_slow_inst_result[26]~q ;
wire \A_wr_data_unfiltered[26]~49_combout ;
wire \A_wr_data_unfiltered[26]~50_combout ;
wire \W_wr_data[26]~q ;
wire \D_src1_reg[26]~20_combout ;
wire \E_src1[26]~q ;
wire \E_alu_result~22_combout ;
wire \D_src2_reg[26]~66_combout ;
wire \D_src2_reg[26]~45_combout ;
wire \D_src2[26]~14_combout ;
wire \D_src2[26]~15_combout ;
wire \E_src2[26]~q ;
wire \Add17~106 ;
wire \Add17~98 ;
wire \Add17~133_sumout ;
wire \D_src2_reg[28]~63_combout ;
wire \D_src2_reg[28]~64_combout ;
wire \D_src2[28]~10_combout ;
wire \D_src2[28]~11_combout ;
wire \E_src2[28]~q ;
wire \E_alu_result~31_combout ;
wire \E_alu_result[28]~combout ;
wire \M_alu_result[28]~q ;
wire \A_inst_result[28]~q ;
wire \M_rot[4]~31_combout ;
wire \A_shift_rot_result~31_combout ;
wire \A_shift_rot_result[28]~q ;
wire \A_slow_inst_result[28]~q ;
wire \A_wr_data_unfiltered[28]~65_combout ;
wire \A_wr_data_unfiltered[28]~66_combout ;
wire \W_wr_data[28]~q ;
wire \D_src1_reg[28]~18_combout ;
wire \E_src1[28]~q ;
wire \E_rot_step1[28]~21_combout ;
wire \M_rot_prestep2[0]~q ;
wire \M_rot[0]~6_combout ;
wire \A_shift_rot_result~6_combout ;
wire \A_shift_rot_result[8]~q ;
wire \A_slow_ld_byte1_data_aligned_nxt[0]~5_combout ;
wire \A_slow_inst_result[8]~q ;
wire \A_wr_data_unfiltered[8]~16_combout ;
wire \A_wr_data_unfiltered[8]~17_combout ;
wire \W_wr_data[8]~q ;
wire \D_src2_reg[8]~13_combout ;
wire \D_src2_reg[8]~97_combout ;
wire \E_logic_result[8]~5_combout ;
wire \E_alu_result[8]~7_combout ;
wire \D_src2_reg[8]~108_combout ;
wire \E_src2[8]~q ;
wire \Add17~1_sumout ;
wire \E_alu_result[8]~combout ;
wire \M_alu_result[8]~q ;
wire \A_inst_result[8]~q ;
wire \A_wr_data_unfiltered[0]~30_combout ;
wire \E_rot_pass0~0_combout ;
wire \M_rot_pass0~q ;
wire \E_rot_sel_fill0~0_combout ;
wire \M_rot_sel_fill0~q ;
wire \M_rot[0]~13_combout ;
wire \A_shift_rot_result~13_combout ;
wire \A_shift_rot_result[0]~q ;
wire \A_wr_data_unfiltered[0]~1_combout ;
wire \A_wr_data_unfiltered[0]~2_combout ;
wire \A_wr_data_unfiltered[0]~31_combout ;
wire \W_wr_data[0]~q ;
wire \D_src1_reg[0]~31_combout ;
wire \E_src1[0]~q ;
wire \Add17~70_cout ;
wire \Add17~58 ;
wire \Add17~54 ;
wire \Add17~26 ;
wire \Add17~30 ;
wire \Add17~34 ;
wire \Add17~17_sumout ;
wire \E_alu_result~10_combout ;
wire \E_alu_result[5]~combout ;
wire \M_alu_result[5]~q ;
wire \A_inst_result[5]~q ;
wire \A_wr_data_unfiltered[5]~22_combout ;
wire \M_rot[5]~9_combout ;
wire \A_shift_rot_result~9_combout ;
wire \A_shift_rot_result[5]~q ;
wire \A_wr_data_unfiltered[5]~23_combout ;
wire \W_wr_data[5]~q ;
wire \D_src1_reg[5]~9_combout ;
wire \E_src1[5]~q ;
wire \E_rot_step1[6]~6_combout ;
wire \M_rot_prestep2[10]~q ;
wire \M_rot[2]~4_combout ;
wire \A_shift_rot_result~4_combout ;
wire \A_shift_rot_result[10]~q ;
wire \A_wr_data_unfiltered[10]~13_combout ;
wire \W_wr_data[10]~q ;
wire \D_src1_reg[10]~4_combout ;
wire \E_src1[10]~q ;
wire \E_rot_step1[10]~7_combout ;
wire \M_rot_prestep2[14]~q ;
wire \M_rot[6]~27_combout ;
wire \A_shift_rot_result~27_combout ;
wire \A_shift_rot_result[14]~q ;
wire \A_slow_ld_byte1_data_aligned_nxt[6]~7_combout ;
wire \A_slow_inst_result[14]~q ;
wire \A_wr_data_unfiltered[14]~58_combout ;
wire \A_wr_data_unfiltered[14]~68_combout ;
wire \W_wr_data[14]~q ;
wire \D_src2_reg[14]~54_combout ;
wire \D_src2_reg[14]~99_combout ;
wire \Add17~125_sumout ;
wire \D_src2_reg[14]~100_combout ;
wire \E_src2[14]~q ;
wire \E_alu_result~27_combout ;
wire \E_alu_result[14]~combout ;
wire \M_alu_result[14]~q ;
wire \A_inst_result[14]~q ;
wire \A_wr_data_unfiltered[6]~20_combout ;
wire \M_rot[6]~8_combout ;
wire \A_shift_rot_result~8_combout ;
wire \A_shift_rot_result[6]~q ;
wire \A_wr_data_unfiltered[6]~21_combout ;
wire \W_wr_data[6]~q ;
wire \D_src1_reg[6]~8_combout ;
wire \E_src1[6]~q ;
wire \Add17~18 ;
wire \Add17~21_sumout ;
wire \E_alu_result~9_combout ;
wire \E_alu_result[6]~combout ;
wire \M_alu_result[6]~q ;
wire \D_src2_reg[6]~16_combout ;
wire \D_src2_reg[6]~17_combout ;
wire \E_src2[6]~q ;
wire \Add17~22 ;
wire \Add17~9_sumout ;
wire \E_alu_result~8_combout ;
wire \E_alu_result[7]~combout ;
wire \M_alu_result[7]~q ;
wire \A_inst_result[7]~q ;
wire \A_wr_data_unfiltered[7]~18_combout ;
wire \M_rot[7]~7_combout ;
wire \A_shift_rot_result~7_combout ;
wire \A_shift_rot_result[7]~q ;
wire \A_wr_data_unfiltered[7]~19_combout ;
wire \W_wr_data[7]~q ;
wire \D_src1_reg[7]~7_combout ;
wire \E_src1[7]~q ;
wire \E_rot_step1[7]~24_combout ;
wire \M_rot_prestep2[11]~q ;
wire \M_rot[3]~3_combout ;
wire \A_shift_rot_result~3_combout ;
wire \A_shift_rot_result[11]~q ;
wire \A_slow_ld_byte1_data_aligned_nxt[3]~2_combout ;
wire \A_slow_inst_result[11]~q ;
wire \A_wr_data_unfiltered[11]~10_combout ;
wire \A_wr_data_unfiltered[11]~11_combout ;
wire \W_wr_data[11]~q ;
wire \D_src2_reg[11]~10_combout ;
wire \D_src2_reg[11]~94_combout ;
wire \E_logic_result[11]~2_combout ;
wire \E_alu_result[11]~4_combout ;
wire \D_src2_reg[11]~120_combout ;
wire \E_src2[11]~q ;
wire \Add17~49_sumout ;
wire \E_alu_result[11]~combout ;
wire \M_alu_result[11]~q ;
wire \A_inst_result[11]~q ;
wire \A_wr_data_unfiltered[3]~26_combout ;
wire \M_rot[3]~11_combout ;
wire \A_shift_rot_result~11_combout ;
wire \A_shift_rot_result[3]~q ;
wire \A_wr_data_unfiltered[3]~27_combout ;
wire \W_wr_data[3]~q ;
wire \D_src1_reg[3]~11_combout ;
wire \E_src1[3]~q ;
wire \Add17~29_sumout ;
wire \E_alu_result~12_combout ;
wire \E_alu_result[3]~combout ;
wire \M_alu_result[3]~q ;
wire \D_src2_reg[3]~22_combout ;
wire \D_src2_reg[3]~23_combout ;
wire \E_src2[3]~q ;
wire \E_rot_pass1~0_combout ;
wire \M_rot_pass1~q ;
wire \M_rot[4]~2_combout ;
wire \A_shift_rot_result~2_combout ;
wire \A_shift_rot_result[12]~q ;
wire \A_slow_ld_byte1_data_aligned_nxt[4]~1_combout ;
wire \A_slow_inst_result[12]~q ;
wire \A_wr_data_unfiltered[12]~8_combout ;
wire \A_wr_data_unfiltered[12]~9_combout ;
wire \W_wr_data[12]~q ;
wire \D_src2_reg[12]~9_combout ;
wire \D_src2_reg[12]~93_combout ;
wire \E_logic_result[12]~1_combout ;
wire \E_alu_result[12]~3_combout ;
wire \D_src2_reg[12]~124_combout ;
wire \E_src2[12]~q ;
wire \Add17~45_sumout ;
wire \E_alu_result[12]~combout ;
wire \M_alu_result[12]~q ;
wire \A_inst_result[12]~q ;
wire \A_wr_data_unfiltered[4]~24_combout ;
wire \M_rot[4]~10_combout ;
wire \A_shift_rot_result~10_combout ;
wire \A_shift_rot_result[4]~q ;
wire \A_wr_data_unfiltered[4]~25_combout ;
wire \W_wr_data[4]~q ;
wire \D_src2_reg[4]~20_combout ;
wire \D_src2_reg[4]~21_combout ;
wire \E_src2[4]~q ;
wire \Add17~33_sumout ;
wire \E_alu_result~11_combout ;
wire \E_alu_result[4]~combout ;
wire \M_alu_result[4]~q ;
wire \A_mem_baddr[4]~q ;
wire \A_dc_fill_has_started_nxt~0_combout ;
wire \A_dc_fill_has_started~q ;
wire \A_dc_fill_starting~0_combout ;
wire \A_dc_fill_dp_offset_nxt[0]~1_combout ;
wire \A_dc_rd_data_cnt[0]~1_combout ;
wire \A_dc_fill_dp_offset[0]~q ;
wire \A_dc_fill_dp_offset_nxt[1]~2_combout ;
wire \A_dc_fill_dp_offset[1]~q ;
wire \A_dc_fill_dp_offset_nxt[2]~0_combout ;
wire \A_dc_fill_dp_offset[2]~q ;
wire \Equal264~0_combout ;
wire \M_ctrl_ld_st_nxt~0_combout ;
wire \M_ctrl_ld_st~q ;
wire \M_valid_mem_d1~0_combout ;
wire \M_valid_mem_d1~q ;
wire \A_mem_baddr[10]~q ;
wire \A_mem_baddr[7]~q ;
wire \A_mem_baddr[6]~q ;
wire \A_mem_baddr[5]~q ;
wire \Equal262~0_combout ;
wire \A_mem_baddr[9]~q ;
wire \A_mem_baddr[8]~q ;
wire \Equal262~1_combout ;
wire \Equal262~2_combout ;
wire \M_A_dc_line_match_d1~q ;
wire \A_dc_fill_need_extra_stall_nxt~combout ;
wire \A_dc_fill_need_extra_stall~q ;
wire \A_dc_rd_data_cnt_nxt[0]~3_combout ;
wire \A_dc_rd_data_cnt[0]~0_combout ;
wire \A_dc_rd_data_cnt[0]~q ;
wire \A_dc_rd_data_cnt_nxt[1]~2_combout ;
wire \A_dc_rd_data_cnt[1]~q ;
wire \A_dc_rd_data_cnt_nxt[2]~1_combout ;
wire \A_dc_rd_data_cnt[2]~q ;
wire \A_dc_rd_data_cnt_nxt[3]~0_combout ;
wire \A_dc_rd_data_cnt[3]~q ;
wire \A_ld_bypass_done~combout ;
wire \A_dc_rd_last_transfer_d1~q ;
wire \A_dc_fill_active_nxt~0_combout ;
wire \A_dc_fill_active~q ;
wire \A_mem_baddr[3]~q ;
wire \A_mem_baddr[2]~q ;
wire \A_dc_fill_wr_data~0_combout ;
wire \A_slow_inst_result_en~0_combout ;
wire \A_slow_inst_result[1]~q ;
wire \A_inst_result[1]~q ;
wire \A_wr_data_unfiltered[1]~28_combout ;
wire \M_rot[1]~12_combout ;
wire \A_shift_rot_result~12_combout ;
wire \A_shift_rot_result[1]~q ;
wire \A_wr_data_unfiltered[1]~29_combout ;
wire \W_wr_data[1]~q ;
wire \D_src2_reg[1]~24_combout ;
wire \D_src2_reg[1]~25_combout ;
wire \E_src2[1]~q ;
wire \Add17~53_sumout ;
wire \E_logic_result[1]~12_combout ;
wire \E_alu_result[1]~combout ;
wire \M_alu_result[1]~q ;
wire \M_ld_align_sh16~0_combout ;
wire \A_ld_align_sh16~q ;
wire \A_slow_ld_byte0_data_aligned_nxt[2]~0_combout ;
wire \A_slow_inst_result[2]~q ;
wire \A_inst_result[2]~q ;
wire \A_wr_data_unfiltered[2]~0_combout ;
wire \M_rot[2]~0_combout ;
wire \A_shift_rot_result~0_combout ;
wire \A_shift_rot_result[2]~q ;
wire \A_wr_data_unfiltered[2]~3_combout ;
wire \W_wr_data[2]~q ;
wire \D_src1_reg[2]~0_combout ;
wire \E_src1[2]~q ;
wire \Add17~25_sumout ;
wire \E_alu_result~1_combout ;
wire \E_alu_result[2]~combout ;
wire \M_alu_result[2]~q ;
wire \D_src2_reg[2]~5_combout ;
wire \D_src2_reg[2]~6_combout ;
wire \E_src2[2]~q ;
wire \E_rot_mask[3]~3_combout ;
wire \M_rot_mask[3]~q ;
wire \M_rot[3]~20_combout ;
wire \A_shift_rot_result~20_combout ;
wire \A_shift_rot_result[27]~q ;
wire \A_slow_inst_result[27]~q ;
wire \A_wr_data_unfiltered[27]~45_combout ;
wire \A_wr_data_unfiltered[27]~46_combout ;
wire \W_wr_data[27]~q ;
wire \D_src1_reg[27]~12_combout ;
wire \E_src1[27]~q ;
wire \Add17~97_sumout ;
wire \D_src2_reg[27]~56_combout ;
wire \D_src2_reg[27]~41_combout ;
wire \D_src2[27]~0_combout ;
wire \D_src2[27]~1_combout ;
wire \E_src2[27]~q ;
wire \E_logic_result[27]~6_combout ;
wire \Equal303~0_combout ;
wire \Equal303~1_combout ;
wire \Equal303~2_combout ;
wire \Equal303~3_combout ;
wire \Equal303~4_combout ;
wire \Equal303~5_combout ;
wire \Equal303~6_combout ;
wire \Equal303~7_combout ;
wire \Equal303~8_combout ;
wire \Equal303~9_combout ;
wire \Equal303~10_combout ;
wire \Equal303~11_combout ;
wire \Equal303~12_combout ;
wire \Equal303~13_combout ;
wire \Equal303~14_combout ;
wire \Equal303~15_combout ;
wire \E_compare_op[1]~q ;
wire \E_br_result~0_combout ;
wire \E_br_result~1_combout ;
wire \E_logic_result[0]~13_combout ;
wire \E_alu_result[0]~13_combout ;
wire \E_alu_result[0]~combout ;
wire \D_src2_reg[0]~26_combout ;
wire \D_src2_reg[0]~27_combout ;
wire \E_src2[0]~q ;
wire \Add17~57_sumout ;
wire \M_data_ram_ld_align_sign_bit_16_hi~0_combout ;
wire \M_data_ram_ld_align_sign_bit_16_hi~q ;
wire \M_data_ram_ld_align_sign_bit~0_combout ;
wire \A_data_ram_ld_align_sign_bit~q ;
wire \M_rot[7]~30_combout ;
wire \A_shift_rot_result~30_combout ;
wire \A_shift_rot_result[31]~q ;
wire \A_slow_inst_result[31]~q ;
wire \A_wr_data_unfiltered[31]~63_combout ;
wire \A_wr_data_unfiltered[31]~64_combout ;
wire \W_wr_data[31]~q ;
wire \D_src1_reg[31]~15_combout ;
wire \E_src1[31]~q ;
wire \Add17~66 ;
wire \Add17~37_sumout ;
wire \D_src2_reg[31]~61_combout ;
wire \D_src2_reg[31]~62_combout ;
wire \D_src2[31]~6_combout ;
wire \D_src2[31]~7_combout ;
wire \E_src2[31]~q ;
wire \Add17~38 ;
wire \Add17~61_sumout ;
wire \E_br_result~2_combout ;
wire \E_ctrl_br_cond~q ;
wire \D_ctrl_flush_pipe_always~0_combout ;
wire \D_ctrl_flush_pipe_always~1_combout ;
wire \E_ctrl_flush_pipe_always~q ;
wire \M_pipe_flush_nxt~0_combout ;
wire \M_pipe_flush~q ;
wire \E_wr_dst_reg_from_D~q ;
wire \E_wr_dst_reg~0_combout ;
wire \E_regnum_b_cmp_F~0_combout ;
wire \E_regnum_b_cmp_F~1_combout ;
wire \E_regnum_b_cmp_F~combout ;
wire \M_regnum_b_cmp_D~q ;
wire \D_data_depend~1_combout ;
wire \D_dep_stall~0_combout ;
wire \F_stall~combout ;
wire \D_iw[5]~q ;
wire \E_iw[5]~q ;
wire \E_ld_st_dcache_management_bus~0_combout ;
wire \M_ctrl_ld_st_bypass_or_dcache_management~q ;
wire \A_mem_stall_nxt~0_combout ;
wire \M_sel_data_master~q ;
wire \M_ctrl_st_nxt~0_combout ;
wire \E_st_cache~0_combout ;
wire \M_ctrl_st_non_bypass~q ;
wire \M_dc_valid_st_cache_hit~0_combout ;
wire \M_dc_potential_hazard_after_st_unfiltered~0_combout ;
wire \M_dc_potential_hazard_after_st_unfiltered~1_combout ;
wire \M_dc_potential_hazard_after_st_unfiltered~2_combout ;
wire \M_dc_potential_hazard_after_st_unfiltered~3_combout ;
wire \M_dc_potential_hazard_after_st_unfiltered~4_combout ;
wire \A_mem_stall_nxt~1_combout ;
wire \E_st_bus~0_combout ;
wire \M_ctrl_st_bypass~q ;
wire \A_ctrl_st_bypass~q ;
wire \M_dc_hit~0_combout ;
wire \M_dc_hit~combout ;
wire \M_dc_valid_st_bypass_hit~0_combout ;
wire \A_dc_valid_st_bypass_hit~q ;
wire \A_st_bypass_transfer_done~combout ;
wire \A_st_bypass_transfer_done_d1~q ;
wire \A_valid~q ;
wire \M_dc_valid_st_cache_hit~1_combout ;
wire \A_dc_valid_st_cache_hit~q ;
wire \M_dc_dirty~combout ;
wire \A_dc_dirty~q ;
wire \Equal193~0_combout ;
wire \M_ctrl_dc_index_wb_inv~q ;
wire \A_ctrl_dc_index_wb_inv~q ;
wire \A_dc_hit~q ;
wire \E_ctrl_dc_addr_inv~0_combout ;
wire \Equal181~0_combout ;
wire \M_ctrl_dc_addr_wb_inv~q ;
wire \A_ctrl_dc_addr_wb_inv~q ;
wire \Equal178~0_combout ;
wire \M_ctrl_dc_nowb_inv~q ;
wire \A_ctrl_dc_nowb_inv~q ;
wire \A_dc_xfer_rd_addr_offset_nxt[0]~1_combout ;
wire \A_dc_xfer_rd_addr_offset[0]~q ;
wire \A_dc_xfer_rd_addr_offset_nxt[1]~0_combout ;
wire \A_dc_xfer_rd_addr_offset[1]~q ;
wire \A_dc_xfer_rd_addr_active_nxt~0_combout ;
wire \A_dc_xfer_rd_addr_active~q ;
wire \A_dc_xfer_rd_addr_offset_nxt[2]~2_combout ;
wire \A_dc_xfer_rd_addr_offset[2]~q ;
wire \A_dc_xfer_rd_addr_done_nxt~combout ;
wire \A_dc_xfer_rd_addr_done~q ;
wire \A_dc_dcache_management_done_nxt~0_combout ;
wire \A_dc_dcache_management_done_nxt~combout ;
wire \A_dc_dcache_management_done~q ;
wire \M_dc_potential_hazard_after_st_unfiltered~5_combout ;
wire \A_dc_potential_hazard_after_st~q ;
wire \A_mem_stall_nxt~2_combout ;
wire \A_mem_stall_nxt~3_combout ;
wire \A_mem_stall_nxt~4_combout ;
wire \A_mem_stall_nxt~5_combout ;
wire \A_mem_stall~q ;
wire \A_stall~combout ;
wire \wait_for_one_post_bret_inst~0_combout ;
wire \wait_for_one_post_bret_inst~q ;
wire \hbreak_req~0_combout ;
wire \latched_oci_tb_hbreak_req_next~0_combout ;
wire \latched_oci_tb_hbreak_req~q ;
wire \F_iw~0_combout ;
wire \F_iw[0]~9_combout ;
wire \D_iw[0]~q ;
wire \Equal171~0_combout ;
wire \D_ctrl_shift_rot~1_combout ;
wire \D_ctrl_late_result~2_combout ;
wire \D_ctrl_late_result~0_combout ;
wire \D_ctrl_late_result~1_combout ;
wire \E_ctrl_late_result~q ;
wire \D_data_depend~0_combout ;
wire \D_valid~combout ;
wire \E_valid_from_D~q ;
wire \E_valid~0_combout ;
wire \E_valid~1_combout ;
wire \M_valid_from_E~q ;
wire \M_dc_want_fill~0_combout ;
wire \E_ld_st_cache~0_combout ;
wire \M_ctrl_ld_st_non_bypass~q ;
wire \M_dc_want_fill~1_combout ;
wire \M_dc_want_fill~combout ;
wire \A_dc_want_fill~q ;
wire \A_dc_xfer_rd_addr_has_started_nxt~0_combout ;
wire \A_dc_xfer_rd_addr_has_started~q ;
wire \A_dc_xfer_rd_addr_starting~0_combout ;
wire \A_dc_xfer_rd_addr_starting~1_combout ;
wire \A_dc_xfer_rd_data_starting~q ;
wire \A_dc_xfer_wr_starting~q ;
wire \A_dc_wb_rd_addr_starting~q ;
wire \A_dc_wb_rd_data_starting~q ;
wire \A_dc_wb_rd_data_first_nxt~0_combout ;
wire \A_dc_wb_rd_data_first~q ;
wire \E_ld_st_bus~0_combout ;
wire \M_ctrl_ld_st_bypass~q ;
wire \A_ctrl_ld_st_bypass~q ;
wire \A_mem_bypass_pending~combout ;
wire \d_address_offset_field[1]~0_combout ;
wire \d_address_offset_field[1]~1_combout ;
wire \d_address_offset_field_nxt[0]~0_combout ;
wire \d_address_offset_field[1]~2_combout ;
wire \d_address_offset_field[1]~3_combout ;
wire \A_st_bypass_delayed~0_combout ;
wire \A_st_bypass_delayed~q ;
wire \A_st_bypass_delayed_started~0_combout ;
wire \A_st_bypass_delayed_started~q ;
wire \d_write_nxt~0_combout ;
wire \d_write_nxt~1_combout ;
wire \A_dc_actual_tag[2]~q ;
wire \A_dc_wb_tag[2]~q ;
wire \A_dc_wb_wr_want_dmaster~combout ;
wire \d_address_tag_field_nxt~0_combout ;
wire \A_mem_baddr[13]~q ;
wire \d_address_tag_field_nxt[2]~1_combout ;
wire \A_dc_actual_tag[1]~q ;
wire \A_dc_wb_tag[1]~q ;
wire \A_mem_baddr[12]~q ;
wire \d_address_tag_field_nxt[1]~2_combout ;
wire \A_dc_actual_tag[0]~q ;
wire \A_dc_wb_tag[0]~q ;
wire \A_mem_baddr[11]~q ;
wire \d_address_tag_field_nxt[0]~3_combout ;
wire \A_dc_wb_line[5]~q ;
wire \d_address_line_field_nxt[5]~0_combout ;
wire \A_dc_wb_line[4]~q ;
wire \d_address_line_field_nxt[4]~1_combout ;
wire \A_dc_wb_line[3]~q ;
wire \d_address_line_field_nxt[3]~2_combout ;
wire \A_dc_wb_line[2]~q ;
wire \d_address_line_field_nxt[2]~3_combout ;
wire \A_dc_wb_line[1]~q ;
wire \d_address_line_field_nxt[1]~4_combout ;
wire \A_dc_wb_line[0]~q ;
wire \d_address_line_field_nxt[0]~5_combout ;
wire \d_address_offset_field_nxt[2]~2_combout ;
wire \d_address_offset_field_nxt[1]~1_combout ;
wire \A_dc_wb_update_av_writedata~combout ;
wire \E_src2_reg[3]~q ;
wire \E_src2_reg[11]~q ;
wire \Equal0~0_combout ;
wire \M_st_data[11]~q ;
wire \A_st_data[11]~q ;
wire \d_writedata_nxt[11]~0_combout ;
wire \d_writedata[14]~0_combout ;
wire \E_mem_byte_en~0_combout ;
wire \M_mem_byte_en[0]~q ;
wire \A_mem_byte_en[0]~q ;
wire \d_byteenable_nxt[1]~0_combout ;
wire \d_byteenable_nxt[0]~1_combout ;
wire \E_src2_reg[2]~q ;
wire \E_src2_reg[10]~q ;
wire \M_st_data[10]~q ;
wire \A_st_data[10]~q ;
wire \d_writedata_nxt[10]~1_combout ;
wire \E_src2_reg[1]~q ;
wire \E_src2_reg[9]~q ;
wire \M_st_data[9]~q ;
wire \A_st_data[9]~q ;
wire \d_writedata_nxt[9]~2_combout ;
wire \E_src2_reg[0]~q ;
wire \E_src2_reg[8]~q ;
wire \M_st_data[8]~q ;
wire \A_st_data[8]~q ;
wire \d_writedata_nxt[8]~3_combout ;
wire \E_src2_reg[5]~q ;
wire \E_src2_reg[13]~q ;
wire \M_st_data[13]~q ;
wire \A_st_data[13]~q ;
wire \d_writedata_nxt[13]~4_combout ;
wire \E_src2_reg[4]~q ;
wire \E_src2_reg[12]~q ;
wire \M_st_data[12]~q ;
wire \A_st_data[12]~q ;
wire \d_writedata_nxt[12]~5_combout ;
wire \D_src2_reg[21]~78_combout ;
wire \D_src2_reg[21]~30_combout ;
wire \E_src2_reg[21]~q ;
wire \M_st_data[21]~q ;
wire \A_st_data[21]~q ;
wire \d_writedata_nxt[21]~6_combout ;
wire \D_src2_reg[20]~79_combout ;
wire \D_src2_reg[20]~32_combout ;
wire \E_src2_reg[20]~q ;
wire \M_st_data[20]~q ;
wire \A_st_data[20]~q ;
wire \d_writedata_nxt[20]~7_combout ;
wire \D_src2_reg[25]~80_combout ;
wire \D_src2_reg[25]~34_combout ;
wire \E_src2_reg[25]~q ;
wire \E_st_data[25]~0_combout ;
wire \M_st_data[25]~q ;
wire \A_st_data[25]~q ;
wire \d_writedata_nxt[25]~8_combout ;
wire \D_src2_reg[17]~36_combout ;
wire \E_src2_reg[17]~q ;
wire \M_st_data[17]~q ;
wire \A_st_data[17]~q ;
wire \d_writedata_nxt[17]~9_combout ;
wire \D_src2_reg[24]~81_combout ;
wire \D_src2_reg[24]~38_combout ;
wire \E_src2_reg[24]~q ;
wire \E_st_data[24]~1_combout ;
wire \M_st_data[24]~q ;
wire \A_st_data[24]~q ;
wire \d_writedata_nxt[24]~10_combout ;
wire \D_src2_reg[16]~40_combout ;
wire \E_src2_reg[16]~q ;
wire \M_st_data[16]~q ;
wire \A_st_data[16]~q ;
wire \d_writedata_nxt[16]~11_combout ;
wire \D_src2_reg[27]~82_combout ;
wire \D_src2_reg[27]~42_combout ;
wire \E_src2_reg[27]~q ;
wire \E_st_data[27]~2_combout ;
wire \M_st_data[27]~q ;
wire \A_st_data[27]~q ;
wire \d_writedata_nxt[27]~12_combout ;
wire \D_src2_reg[19]~83_combout ;
wire \D_src2_reg[19]~44_combout ;
wire \E_src2_reg[19]~q ;
wire \M_st_data[19]~q ;
wire \A_st_data[19]~q ;
wire \d_writedata_nxt[19]~13_combout ;
wire \D_src2_reg[26]~84_combout ;
wire \D_src2_reg[26]~46_combout ;
wire \E_src2_reg[26]~q ;
wire \E_st_data[26]~3_combout ;
wire \M_st_data[26]~q ;
wire \A_st_data[26]~q ;
wire \d_writedata_nxt[26]~14_combout ;
wire \D_src2_reg[18]~85_combout ;
wire \D_src2_reg[18]~48_combout ;
wire \E_src2_reg[18]~q ;
wire \M_st_data[18]~q ;
wire \A_st_data[18]~q ;
wire \d_writedata_nxt[18]~15_combout ;
wire \E_src2_reg[7]~q ;
wire \D_src2_reg[23]~86_combout ;
wire \D_src2_reg[23]~50_combout ;
wire \E_src2_reg[23]~q ;
wire \M_st_data[23]~q ;
wire \A_st_data[23]~q ;
wire \d_writedata_nxt[23]~16_combout ;
wire \E_src2_reg[15]~q ;
wire \M_st_data[15]~q ;
wire \A_st_data[15]~q ;
wire \d_writedata_nxt[15]~17_combout ;
wire \E_src2_reg[6]~q ;
wire \D_src2_reg[22]~87_combout ;
wire \D_src2_reg[22]~53_combout ;
wire \E_src2_reg[22]~q ;
wire \M_st_data[22]~q ;
wire \A_st_data[22]~q ;
wire \d_writedata_nxt[22]~18_combout ;
wire \E_src2_reg[14]~q ;
wire \M_st_data[14]~q ;
wire \A_st_data[14]~q ;
wire \d_writedata_nxt[14]~19_combout ;
wire \A_ld_bypass_delayed~0_combout ;
wire \A_ld_bypass_delayed~q ;
wire \A_ld_bypass_delayed_started~0_combout ;
wire \A_ld_bypass_delayed_started~q ;
wire \d_read_nxt~0_combout ;
wire \d_read_nxt~1_combout ;
wire \A_dc_rd_addr_cnt_nxt[0]~3_combout ;
wire \A_dc_rd_addr_cnt[1]~0_combout ;
wire \A_dc_rd_addr_cnt[0]~q ;
wire \A_dc_rd_addr_cnt_nxt[1]~2_combout ;
wire \A_dc_rd_addr_cnt[1]~q ;
wire \A_dc_rd_addr_cnt_nxt[2]~1_combout ;
wire \A_dc_rd_addr_cnt[2]~q ;
wire \Add15~0_combout ;
wire \A_dc_rd_addr_cnt_nxt[3]~0_combout ;
wire \A_dc_rd_addr_cnt[3]~q ;
wire \d_read_nxt~2_combout ;
wire \E_mem_byte_en[1]~1_combout ;
wire \M_mem_byte_en[1]~q ;
wire \A_mem_byte_en[1]~q ;
wire \d_byteenable_nxt[1]~2_combout ;
wire \M_st_data[2]~q ;
wire \A_st_data[2]~q ;
wire \d_writedata_nxt[2]~20_combout ;
wire \M_st_data[0]~q ;
wire \A_st_data[0]~q ;
wire \d_writedata_nxt[0]~21_combout ;
wire \M_st_data[3]~q ;
wire \A_st_data[3]~q ;
wire \d_writedata_nxt[3]~22_combout ;
wire \M_st_data[1]~q ;
wire \A_st_data[1]~q ;
wire \d_writedata_nxt[1]~23_combout ;
wire \hbreak_enabled~0_combout ;
wire \F_ic_fill_same_tag_line~0_combout ;
wire \F_ic_fill_same_tag_line~1_combout ;
wire \F_ic_fill_same_tag_line~2_combout ;
wire \F_ic_fill_same_tag_line~3_combout ;
wire \F_ic_fill_same_tag_line~combout ;
wire \D_ic_fill_same_tag_line~q ;
wire \E_ctrl_invalidate_i~0_combout ;
wire \E_ctrl_invalidate_i~1_combout ;
wire \M_ctrl_invalidate_i~q ;
wire \ic_tag_clr_valid_bits_nxt~0_combout ;
wire \ic_fill_prevent_refill_nxt~combout ;
wire \ic_fill_prevent_refill~q ;
wire \D_ic_fill_starting~0_combout ;
wire \ic_fill_initial_offset[2]~q ;
wire \D_ic_fill_starting_d1~q ;
wire \ic_fill_initial_offset[0]~q ;
wire \ic_fill_dp_offset_nxt[0]~1_combout ;
wire \i_readdatavalid_d1~q ;
wire \ic_fill_dp_offset_en~0_combout ;
wire \ic_fill_dp_offset[0]~q ;
wire \ic_fill_initial_offset[1]~q ;
wire \ic_fill_dp_offset_nxt[1]~2_combout ;
wire \ic_fill_dp_offset[1]~q ;
wire \ic_fill_dp_offset[2]~q ;
wire \ic_fill_dp_offset_nxt[2]~0_combout ;
wire \ic_fill_active_nxt~0_combout ;
wire \ic_fill_active_nxt~1_combout ;
wire \ic_fill_active~q ;
wire \ic_fill_ap_cnt_nxt[0]~3_combout ;
wire \ic_fill_ap_cnt[1]~0_combout ;
wire \ic_fill_ap_cnt[0]~q ;
wire \ic_fill_ap_cnt_nxt[1]~2_combout ;
wire \ic_fill_ap_cnt[1]~q ;
wire \ic_fill_ap_cnt_nxt[2]~1_combout ;
wire \ic_fill_ap_cnt[2]~q ;
wire \ic_fill_ap_cnt_nxt[3]~0_combout ;
wire \ic_fill_ap_cnt[3]~q ;
wire \i_read_nxt~0_combout ;
wire \i_read_nxt~1_combout ;
wire \ic_tag_wraddress_nxt~0_combout ;
wire \M_st_data[6]~q ;
wire \A_st_data[6]~q ;
wire \d_writedata_nxt[6]~24_combout ;
wire \M_st_data[4]~q ;
wire \A_st_data[4]~q ;
wire \d_writedata_nxt[4]~25_combout ;
wire \M_st_data[7]~q ;
wire \A_st_data[7]~q ;
wire \d_writedata_nxt[7]~26_combout ;
wire \M_st_data[5]~q ;
wire \A_st_data[5]~q ;
wire \d_writedata_nxt[5]~27_combout ;
wire \ic_tag_wraddress_nxt~1_combout ;
wire \ic_fill_ap_offset_nxt[0]~0_combout ;
wire \ic_tag_wraddress_nxt~2_combout ;
wire \ic_tag_wraddress_nxt~3_combout ;
wire \ic_fill_ap_offset_nxt[2]~1_combout ;
wire \ic_fill_ap_offset_nxt[1]~2_combout ;
wire \ic_tag_wraddress_nxt~4_combout ;
wire \ic_tag_wraddress_nxt~5_combout ;
wire \ic_tag_wraddress_nxt~6_combout ;
wire \E_mem_byte_en[2]~2_combout ;
wire \M_mem_byte_en[2]~q ;
wire \A_mem_byte_en[2]~q ;
wire \d_byteenable_nxt[2]~3_combout ;
wire \E_mem_byte_en[3]~3_combout ;
wire \M_mem_byte_en[3]~q ;
wire \A_mem_byte_en[3]~q ;
wire \d_byteenable_nxt[3]~4_combout ;
wire \D_src2_reg[31]~90_combout ;
wire \D_src2_reg[31]~75_combout ;
wire \E_src2_reg[31]~q ;
wire \E_st_data[31]~5_combout ;
wire \M_st_data[31]~q ;
wire \A_st_data[31]~q ;
wire \d_writedata_nxt[31]~28_combout ;
wire \D_src2_reg[29]~88_combout ;
wire \D_src2_reg[29]~74_combout ;
wire \E_src2_reg[29]~q ;
wire \E_st_data[29]~4_combout ;
wire \M_st_data[29]~q ;
wire \A_st_data[29]~q ;
wire \d_writedata_nxt[29]~29_combout ;
wire \D_src2_reg[28]~91_combout ;
wire \D_src2_reg[28]~76_combout ;
wire \E_src2_reg[28]~q ;
wire \E_st_data[28]~6_combout ;
wire \M_st_data[28]~q ;
wire \A_st_data[28]~q ;
wire \d_writedata_nxt[28]~30_combout ;
wire \D_src2_reg[30]~89_combout ;
wire \D_src2_reg[30]~77_combout ;
wire \E_src2_reg[30]~q ;
wire \E_st_data[30]~7_combout ;
wire \M_st_data[30]~q ;
wire \A_st_data[30]~q ;
wire \d_writedata_nxt[30]~31_combout ;


embedded_system_embedded_system_nios2_qsys_0_mult_cell the_embedded_system_nios2_qsys_0_mult_cell(
	.Add0(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~1_sumout ),
	.Add01(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~5_sumout ),
	.Add02(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~9_sumout ),
	.Add03(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~13_sumout ),
	.Add04(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~17_sumout ),
	.Add05(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~21_sumout ),
	.Add06(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~25_sumout ),
	.Add07(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~29_sumout ),
	.Add08(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~33_sumout ),
	.Add09(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~37_sumout ),
	.Add010(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~41_sumout ),
	.Add011(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~45_sumout ),
	.Add012(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~49_sumout ),
	.Add013(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~53_sumout ),
	.Add014(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~57_sumout ),
	.Add015(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~61_sumout ),
	.A_mul_src2_0(\A_mul_src2[0]~q ),
	.A_mul_src2_1(\A_mul_src2[1]~q ),
	.A_mul_src2_2(\A_mul_src2[2]~q ),
	.A_mul_src2_3(\A_mul_src2[3]~q ),
	.A_mul_src2_4(\A_mul_src2[4]~q ),
	.A_mul_src2_5(\A_mul_src2[5]~q ),
	.A_mul_src2_6(\A_mul_src2[6]~q ),
	.A_mul_src2_7(\A_mul_src2[7]~q ),
	.A_mul_src2_8(\A_mul_src2[8]~q ),
	.A_mul_src2_9(\A_mul_src2[9]~q ),
	.A_mul_src2_10(\A_mul_src2[10]~q ),
	.A_mul_src2_11(\A_mul_src2[11]~q ),
	.A_mul_src2_12(\A_mul_src2[12]~q ),
	.A_mul_src2_13(\A_mul_src2[13]~q ),
	.A_mul_src2_14(\A_mul_src2[14]~q ),
	.A_mul_src2_15(\A_mul_src2[15]~q ),
	.A_mul_src1_0(\A_mul_src1[0]~q ),
	.A_mul_src1_1(\A_mul_src1[1]~q ),
	.A_mul_src1_2(\A_mul_src1[2]~q ),
	.A_mul_src1_3(\A_mul_src1[3]~q ),
	.A_mul_src1_4(\A_mul_src1[4]~q ),
	.A_mul_src1_5(\A_mul_src1[5]~q ),
	.A_mul_src1_6(\A_mul_src1[6]~q ),
	.A_mul_src1_7(\A_mul_src1[7]~q ),
	.A_mul_src1_8(\A_mul_src1[8]~q ),
	.A_mul_src1_9(\A_mul_src1[9]~q ),
	.A_mul_src1_10(\A_mul_src1[10]~q ),
	.A_mul_src1_11(\A_mul_src1[11]~q ),
	.A_mul_src1_12(\A_mul_src1[12]~q ),
	.A_mul_src1_13(\A_mul_src1[13]~q ),
	.A_mul_src1_14(\A_mul_src1[14]~q ),
	.A_mul_src1_15(\A_mul_src1[15]~q ),
	.A_mul_src1_16(\A_mul_src1[16]~q ),
	.A_mul_src1_17(\A_mul_src1[17]~q ),
	.A_mul_src1_18(\A_mul_src1[18]~q ),
	.A_mul_src1_19(\A_mul_src1[19]~q ),
	.A_mul_src1_20(\A_mul_src1[20]~q ),
	.A_mul_src1_21(\A_mul_src1[21]~q ),
	.A_mul_src1_22(\A_mul_src1[22]~q ),
	.A_mul_src1_23(\A_mul_src1[23]~q ),
	.A_mul_src1_24(\A_mul_src1[24]~q ),
	.A_mul_src1_25(\A_mul_src1[25]~q ),
	.A_mul_src1_26(\A_mul_src1[26]~q ),
	.A_mul_src1_27(\A_mul_src1[27]~q ),
	.A_mul_src1_28(\A_mul_src1[28]~q ),
	.A_mul_src1_29(\A_mul_src1[29]~q ),
	.A_mul_src1_30(\A_mul_src1[30]~q ),
	.A_mul_src1_31(\A_mul_src1[31]~q ),
	.hq3myc14108phmpo7y7qmhbp98hy0vq(\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.data_out_wire_2(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.data_out_wire_13(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.data_out_wire_12(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.data_out_wire_11(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.data_out_wire_10(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.data_out_wire_9(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.data_out_wire_8(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.data_out_wire_7(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.data_out_wire_6(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.data_out_wire_5(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.data_out_wire_4(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.data_out_wire_3(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.data_out_wire_1(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.data_out_wire_0(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.data_out_wire_15(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.data_out_wire_14(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_dc_victim_module embedded_system_nios2_qsys_0_dc_victim(
	.q_b_11(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_13(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_21(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_25(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_17(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_24(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_16(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_27(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_19(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_26(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_18(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_23(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_15(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_22(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_14(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[14] ),
	.A_dc_xfer_wr_data_11(\A_dc_xfer_wr_data[11]~q ),
	.A_dc_xfer_wr_data_10(\A_dc_xfer_wr_data[10]~q ),
	.A_dc_xfer_wr_data_9(\A_dc_xfer_wr_data[9]~q ),
	.A_dc_xfer_wr_data_8(\A_dc_xfer_wr_data[8]~q ),
	.A_dc_xfer_wr_data_13(\A_dc_xfer_wr_data[13]~q ),
	.A_dc_xfer_wr_data_12(\A_dc_xfer_wr_data[12]~q ),
	.q_b_2(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_0(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_3(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_1(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[1] ),
	.A_dc_xfer_wr_data_21(\A_dc_xfer_wr_data[21]~q ),
	.A_dc_xfer_wr_data_20(\A_dc_xfer_wr_data[20]~q ),
	.A_dc_xfer_wr_data_25(\A_dc_xfer_wr_data[25]~q ),
	.A_dc_xfer_wr_data_17(\A_dc_xfer_wr_data[17]~q ),
	.A_dc_xfer_wr_data_24(\A_dc_xfer_wr_data[24]~q ),
	.A_dc_xfer_wr_data_16(\A_dc_xfer_wr_data[16]~q ),
	.A_dc_xfer_wr_data_27(\A_dc_xfer_wr_data[27]~q ),
	.A_dc_xfer_wr_data_19(\A_dc_xfer_wr_data[19]~q ),
	.A_dc_xfer_wr_data_26(\A_dc_xfer_wr_data[26]~q ),
	.A_dc_xfer_wr_data_18(\A_dc_xfer_wr_data[18]~q ),
	.A_dc_xfer_wr_data_23(\A_dc_xfer_wr_data[23]~q ),
	.A_dc_xfer_wr_data_15(\A_dc_xfer_wr_data[15]~q ),
	.A_dc_xfer_wr_data_22(\A_dc_xfer_wr_data[22]~q ),
	.A_dc_xfer_wr_data_14(\A_dc_xfer_wr_data[14]~q ),
	.A_dc_xfer_wr_data_2(\A_dc_xfer_wr_data[2]~q ),
	.A_dc_xfer_wr_data_0(\A_dc_xfer_wr_data[0]~q ),
	.A_dc_xfer_wr_data_3(\A_dc_xfer_wr_data[3]~q ),
	.q_b_6(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_4(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_7(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_5(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[5] ),
	.A_dc_xfer_wr_data_1(\A_dc_xfer_wr_data[1]~q ),
	.A_dc_xfer_wr_data_6(\A_dc_xfer_wr_data[6]~q ),
	.A_dc_xfer_wr_data_4(\A_dc_xfer_wr_data[4]~q ),
	.A_dc_xfer_wr_data_7(\A_dc_xfer_wr_data[7]~q ),
	.A_dc_xfer_wr_data_5(\A_dc_xfer_wr_data[5]~q ),
	.q_b_31(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_29(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_28(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_30(\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[30] ),
	.A_dc_xfer_wr_data_31(\A_dc_xfer_wr_data[31]~q ),
	.A_dc_xfer_wr_data_29(\A_dc_xfer_wr_data[29]~q ),
	.A_dc_xfer_wr_data_28(\A_dc_xfer_wr_data[28]~q ),
	.A_dc_xfer_wr_data_30(\A_dc_xfer_wr_data[30]~q ),
	.A_dc_xfer_wr_active(\A_dc_xfer_wr_active~q ),
	.A_dc_wb_rd_en(\A_dc_wb_rd_en~combout ),
	.A_dc_xfer_wr_offset_0(\A_dc_xfer_wr_offset[0]~q ),
	.A_dc_xfer_wr_offset_1(\A_dc_xfer_wr_offset[1]~q ),
	.A_dc_xfer_wr_offset_2(\A_dc_xfer_wr_offset[2]~q ),
	.A_dc_wb_rd_addr_offset_0(\A_dc_wb_rd_addr_offset[0]~q ),
	.A_dc_wb_rd_addr_offset_1(\A_dc_wb_rd_addr_offset[1]~q ),
	.A_dc_wb_rd_addr_offset_2(\A_dc_wb_rd_addr_offset[2]~q ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_dc_data_module embedded_system_nios2_qsys_0_dc_data(
	.q_b_11(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_13(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_21(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_25(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_17(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_24(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_16(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_27(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_19(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_26(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_18(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_23(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_15(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_22(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_14(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_2(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_29(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_7(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_31(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_28(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_6(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_30(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_5(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_3(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_1(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ),
	.dc_data_wr_port_en(\dc_data_wr_port_en~combout ),
	.dc_data_wr_port_data_11(\dc_data_wr_port_data[11]~1_combout ),
	.dc_data_wr_port_addr_0(\dc_data_wr_port_addr[0]~0_combout ),
	.dc_data_wr_port_addr_1(\dc_data_wr_port_addr[1]~1_combout ),
	.dc_data_wr_port_addr_2(\dc_data_wr_port_addr[2]~2_combout ),
	.dc_data_wr_port_addr_3(\dc_data_wr_port_addr[3]~3_combout ),
	.dc_data_wr_port_addr_4(\dc_data_wr_port_addr[4]~4_combout ),
	.dc_data_wr_port_addr_5(\dc_data_wr_port_addr[5]~5_combout ),
	.dc_data_wr_port_addr_6(\dc_data_wr_port_addr[6]~6_combout ),
	.dc_data_wr_port_addr_7(\dc_data_wr_port_addr[7]~7_combout ),
	.dc_data_wr_port_addr_8(\dc_data_wr_port_addr[8]~8_combout ),
	.dc_data_rd_port_addr_0(\dc_data_rd_port_addr[0]~0_combout ),
	.dc_data_rd_port_addr_1(\dc_data_rd_port_addr[1]~1_combout ),
	.dc_data_rd_port_addr_2(\dc_data_rd_port_addr[2]~2_combout ),
	.dc_data_rd_port_addr_3(\dc_data_rd_port_addr[3]~3_combout ),
	.dc_data_rd_port_addr_4(\dc_data_rd_port_addr[4]~4_combout ),
	.dc_data_rd_port_addr_5(\dc_data_rd_port_addr[5]~5_combout ),
	.dc_data_rd_port_addr_6(\dc_data_rd_port_addr[6]~6_combout ),
	.dc_data_rd_port_addr_7(\dc_data_rd_port_addr[7]~7_combout ),
	.dc_data_rd_port_addr_8(\dc_data_rd_port_addr[8]~8_combout ),
	.dc_data_wr_port_data_10(\dc_data_wr_port_data[10]~2_combout ),
	.dc_data_wr_port_data_9(\dc_data_wr_port_data[9]~3_combout ),
	.dc_data_wr_port_data_8(\dc_data_wr_port_data[8]~4_combout ),
	.dc_data_wr_port_data_13(\dc_data_wr_port_data[13]~5_combout ),
	.dc_data_wr_port_data_12(\dc_data_wr_port_data[12]~6_combout ),
	.dc_data_wr_port_data_21(\dc_data_wr_port_data[21]~8_combout ),
	.dc_data_wr_port_data_20(\dc_data_wr_port_data[20]~9_combout ),
	.dc_data_wr_port_data_25(\dc_data_wr_port_data[25]~11_combout ),
	.dc_data_wr_port_data_17(\dc_data_wr_port_data[17]~12_combout ),
	.dc_data_wr_port_data_24(\dc_data_wr_port_data[24]~13_combout ),
	.dc_data_wr_port_data_16(\dc_data_wr_port_data[16]~14_combout ),
	.dc_data_wr_port_data_27(\dc_data_wr_port_data[27]~15_combout ),
	.dc_data_wr_port_data_19(\dc_data_wr_port_data[19]~16_combout ),
	.dc_data_wr_port_data_26(\dc_data_wr_port_data[26]~17_combout ),
	.dc_data_wr_port_data_18(\dc_data_wr_port_data[18]~18_combout ),
	.dc_data_wr_port_data_23(\dc_data_wr_port_data[23]~19_combout ),
	.dc_data_wr_port_data_15(\dc_data_wr_port_data[15]~20_combout ),
	.dc_data_wr_port_data_22(\dc_data_wr_port_data[22]~21_combout ),
	.dc_data_wr_port_data_14(\dc_data_wr_port_data[14]~22_combout ),
	.dc_data_wr_port_data_2(\dc_data_wr_port_data[2]~24_combout ),
	.dc_data_wr_port_data_29(\dc_data_wr_port_data[29]~25_combout ),
	.dc_data_wr_port_data_7(\dc_data_wr_port_data[7]~26_combout ),
	.dc_data_wr_port_data_31(\dc_data_wr_port_data[31]~27_combout ),
	.dc_data_wr_port_data_28(\dc_data_wr_port_data[28]~28_combout ),
	.dc_data_wr_port_data_6(\dc_data_wr_port_data[6]~29_combout ),
	.dc_data_wr_port_data_30(\dc_data_wr_port_data[30]~30_combout ),
	.dc_data_wr_port_data_5(\dc_data_wr_port_data[5]~31_combout ),
	.dc_data_wr_port_data_4(\dc_data_wr_port_data[4]~32_combout ),
	.dc_data_wr_port_data_3(\dc_data_wr_port_data[3]~33_combout ),
	.dc_data_wr_port_data_1(\dc_data_wr_port_data[1]~34_combout ),
	.dc_data_wr_port_data_0(\dc_data_wr_port_data[0]~35_combout ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_dc_tag_module embedded_system_nios2_qsys_0_dc_tag(
	.q_b_1(\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_2(\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_3(\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_0(\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_4(\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[4] ),
	.dc_tag_wr_port_en(\dc_tag_wr_port_en~combout ),
	.dc_tag_wr_port_data_1(\dc_tag_wr_port_data[1]~0_combout ),
	.dc_tag_wr_port_addr_0(\dc_tag_wr_port_addr[0]~1_combout ),
	.dc_tag_wr_port_addr_1(\dc_tag_wr_port_addr[1]~2_combout ),
	.dc_tag_wr_port_addr_2(\dc_tag_wr_port_addr[2]~3_combout ),
	.dc_tag_wr_port_addr_3(\dc_tag_wr_port_addr[3]~4_combout ),
	.dc_tag_wr_port_addr_4(\dc_tag_wr_port_addr[4]~5_combout ),
	.dc_tag_wr_port_addr_5(\dc_tag_wr_port_addr[5]~6_combout ),
	.dc_tag_rd_port_addr_0(\dc_tag_rd_port_addr[0]~0_combout ),
	.dc_tag_rd_port_addr_1(\dc_tag_rd_port_addr[1]~1_combout ),
	.dc_tag_rd_port_addr_2(\dc_tag_rd_port_addr[2]~2_combout ),
	.dc_tag_rd_port_addr_3(\dc_tag_rd_port_addr[3]~3_combout ),
	.dc_tag_rd_port_addr_4(\dc_tag_rd_port_addr[4]~4_combout ),
	.dc_tag_rd_port_addr_5(\dc_tag_rd_port_addr[5]~5_combout ),
	.dc_tag_wr_port_data_2(\dc_tag_wr_port_data[2]~1_combout ),
	.dc_tag_wr_port_data_3(\dc_tag_wr_port_data[3]~2_combout ),
	.dc_tag_wr_port_data_0(\dc_tag_wr_port_data[0]~3_combout ),
	.dc_tag_wr_port_data_4(\dc_tag_wr_port_data[4]~4_combout ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_register_bank_b_module embedded_system_nios2_qsys_0_register_bank_b(
	.q_b_2(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_13(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_5(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_3(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_1(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_21(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_25(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_17(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_24(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_16(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_27(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_19(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_26(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_18(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_23(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_15(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_22(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_14(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_29(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_30(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_31(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_28(\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.A_wr_data_unfiltered_2(\A_wr_data_unfiltered[2]~3_combout ),
	.A_wr_data_unfiltered_13(\A_wr_data_unfiltered[13]~7_combout ),
	.A_wr_data_unfiltered_12(\A_wr_data_unfiltered[12]~9_combout ),
	.A_wr_data_unfiltered_11(\A_wr_data_unfiltered[11]~11_combout ),
	.A_wr_data_unfiltered_10(\A_wr_data_unfiltered[10]~13_combout ),
	.A_wr_data_unfiltered_9(\A_wr_data_unfiltered[9]~15_combout ),
	.A_wr_data_unfiltered_8(\A_wr_data_unfiltered[8]~17_combout ),
	.A_wr_data_unfiltered_7(\A_wr_data_unfiltered[7]~19_combout ),
	.A_wr_data_unfiltered_6(\A_wr_data_unfiltered[6]~21_combout ),
	.A_wr_data_unfiltered_5(\A_wr_data_unfiltered[5]~23_combout ),
	.A_wr_data_unfiltered_4(\A_wr_data_unfiltered[4]~25_combout ),
	.A_wr_data_unfiltered_3(\A_wr_data_unfiltered[3]~27_combout ),
	.A_wr_data_unfiltered_1(\A_wr_data_unfiltered[1]~29_combout ),
	.A_wr_data_unfiltered_0(\A_wr_data_unfiltered[0]~31_combout ),
	.A_wr_data_unfiltered_21(\A_wr_data_unfiltered[21]~34_combout ),
	.A_wr_data_unfiltered_20(\A_wr_data_unfiltered[20]~36_combout ),
	.A_wr_data_unfiltered_25(\A_wr_data_unfiltered[25]~38_combout ),
	.A_wr_data_unfiltered_17(\A_wr_data_unfiltered[17]~40_combout ),
	.A_wr_data_unfiltered_24(\A_wr_data_unfiltered[24]~42_combout ),
	.A_wr_data_unfiltered_16(\A_wr_data_unfiltered[16]~44_combout ),
	.A_wr_data_unfiltered_27(\A_wr_data_unfiltered[27]~46_combout ),
	.A_wr_data_unfiltered_19(\A_wr_data_unfiltered[19]~48_combout ),
	.A_wr_data_unfiltered_26(\A_wr_data_unfiltered[26]~50_combout ),
	.A_wr_data_unfiltered_18(\A_wr_data_unfiltered[18]~52_combout ),
	.A_wr_data_unfiltered_23(\A_wr_data_unfiltered[23]~54_combout ),
	.A_wr_data_unfiltered_22(\A_wr_data_unfiltered[22]~57_combout ),
	.A_wr_data_unfiltered_29(\A_wr_data_unfiltered[29]~60_combout ),
	.A_wr_data_unfiltered_30(\A_wr_data_unfiltered[30]~62_combout ),
	.A_wr_data_unfiltered_31(\A_wr_data_unfiltered[31]~64_combout ),
	.A_wr_data_unfiltered_28(\A_wr_data_unfiltered[28]~66_combout ),
	.A_wr_data_unfiltered_15(\A_wr_data_unfiltered[15]~67_combout ),
	.A_wr_data_unfiltered_14(\A_wr_data_unfiltered[14]~68_combout ),
	.A_dst_regnum_from_M_4(\A_dst_regnum_from_M[4]~q ),
	.A_wr_dst_reg_from_M(\A_wr_dst_reg_from_M~q ),
	.A_dst_regnum_from_M_0(\A_dst_regnum_from_M[0]~q ),
	.A_dst_regnum_from_M_1(\A_dst_regnum_from_M[1]~q ),
	.A_dst_regnum_from_M_2(\A_dst_regnum_from_M[2]~q ),
	.A_dst_regnum_from_M_3(\A_dst_regnum_from_M[3]~q ),
	.rf_b_rd_port_addr_0(\rf_b_rd_port_addr[0]~0_combout ),
	.rf_b_rd_port_addr_1(\rf_b_rd_port_addr[1]~1_combout ),
	.rf_b_rd_port_addr_2(\rf_b_rd_port_addr[2]~2_combout ),
	.rf_b_rd_port_addr_3(\rf_b_rd_port_addr[3]~3_combout ),
	.rf_b_rd_port_addr_4(\rf_b_rd_port_addr[4]~4_combout ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_register_bank_a_module embedded_system_nios2_qsys_0_register_bank_a(
	.q_b_2(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_13(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_12(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_10(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_8(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_7(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_5(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_4(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_3(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_27(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_29(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_30(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_31(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_17(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_16(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_28(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_18(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_26(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_19(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_21(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_15(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_25(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_20(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_22(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_14(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_24(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_23(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_1(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.A_wr_data_unfiltered_2(\A_wr_data_unfiltered[2]~3_combout ),
	.A_wr_data_unfiltered_13(\A_wr_data_unfiltered[13]~7_combout ),
	.A_wr_data_unfiltered_12(\A_wr_data_unfiltered[12]~9_combout ),
	.A_wr_data_unfiltered_11(\A_wr_data_unfiltered[11]~11_combout ),
	.A_wr_data_unfiltered_10(\A_wr_data_unfiltered[10]~13_combout ),
	.A_wr_data_unfiltered_9(\A_wr_data_unfiltered[9]~15_combout ),
	.A_wr_data_unfiltered_8(\A_wr_data_unfiltered[8]~17_combout ),
	.A_wr_data_unfiltered_7(\A_wr_data_unfiltered[7]~19_combout ),
	.A_wr_data_unfiltered_6(\A_wr_data_unfiltered[6]~21_combout ),
	.A_wr_data_unfiltered_5(\A_wr_data_unfiltered[5]~23_combout ),
	.A_wr_data_unfiltered_4(\A_wr_data_unfiltered[4]~25_combout ),
	.A_wr_data_unfiltered_3(\A_wr_data_unfiltered[3]~27_combout ),
	.A_wr_data_unfiltered_1(\A_wr_data_unfiltered[1]~29_combout ),
	.A_wr_data_unfiltered_0(\A_wr_data_unfiltered[0]~31_combout ),
	.A_wr_data_unfiltered_21(\A_wr_data_unfiltered[21]~34_combout ),
	.A_wr_data_unfiltered_20(\A_wr_data_unfiltered[20]~36_combout ),
	.A_wr_data_unfiltered_25(\A_wr_data_unfiltered[25]~38_combout ),
	.A_wr_data_unfiltered_17(\A_wr_data_unfiltered[17]~40_combout ),
	.A_wr_data_unfiltered_24(\A_wr_data_unfiltered[24]~42_combout ),
	.A_wr_data_unfiltered_16(\A_wr_data_unfiltered[16]~44_combout ),
	.A_wr_data_unfiltered_27(\A_wr_data_unfiltered[27]~46_combout ),
	.A_wr_data_unfiltered_19(\A_wr_data_unfiltered[19]~48_combout ),
	.A_wr_data_unfiltered_26(\A_wr_data_unfiltered[26]~50_combout ),
	.A_wr_data_unfiltered_18(\A_wr_data_unfiltered[18]~52_combout ),
	.A_wr_data_unfiltered_23(\A_wr_data_unfiltered[23]~54_combout ),
	.A_wr_data_unfiltered_22(\A_wr_data_unfiltered[22]~57_combout ),
	.A_wr_data_unfiltered_29(\A_wr_data_unfiltered[29]~60_combout ),
	.A_wr_data_unfiltered_30(\A_wr_data_unfiltered[30]~62_combout ),
	.A_wr_data_unfiltered_31(\A_wr_data_unfiltered[31]~64_combout ),
	.A_wr_data_unfiltered_28(\A_wr_data_unfiltered[28]~66_combout ),
	.A_wr_data_unfiltered_15(\A_wr_data_unfiltered[15]~67_combout ),
	.A_wr_data_unfiltered_14(\A_wr_data_unfiltered[14]~68_combout ),
	.A_dst_regnum_from_M_4(\A_dst_regnum_from_M[4]~q ),
	.A_wr_dst_reg_from_M(\A_wr_dst_reg_from_M~q ),
	.A_dst_regnum_from_M_0(\A_dst_regnum_from_M[0]~q ),
	.A_dst_regnum_from_M_1(\A_dst_regnum_from_M[1]~q ),
	.A_dst_regnum_from_M_2(\A_dst_regnum_from_M[2]~q ),
	.A_dst_regnum_from_M_3(\A_dst_regnum_from_M[3]~q ),
	.rf_a_rd_port_addr_0(\rf_a_rd_port_addr[0]~0_combout ),
	.rf_a_rd_port_addr_1(\rf_a_rd_port_addr[1]~1_combout ),
	.rf_a_rd_port_addr_2(\rf_a_rd_port_addr[2]~2_combout ),
	.rf_a_rd_port_addr_3(\rf_a_rd_port_addr[3]~3_combout ),
	.rf_a_rd_port_addr_4(\rf_a_rd_port_addr[4]~4_combout ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_bht_module embedded_system_nios2_qsys_0_bht(
	.q_b_1(\embedded_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_0(\embedded_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[0] ),
	.F_stall(\F_stall~combout ),
	.M_bht_wr_en_unfiltered(\M_bht_wr_en_unfiltered~combout ),
	.M_bht_wr_data_unfiltered_1(\M_bht_wr_data_unfiltered[1]~0_combout ),
	.M_bht_ptr_unfiltered_0(\M_bht_ptr_unfiltered[0]~q ),
	.M_bht_ptr_unfiltered_1(\M_bht_ptr_unfiltered[1]~q ),
	.M_bht_ptr_unfiltered_2(\M_bht_ptr_unfiltered[2]~q ),
	.M_bht_ptr_unfiltered_3(\M_bht_ptr_unfiltered[3]~q ),
	.M_bht_ptr_unfiltered_4(\M_bht_ptr_unfiltered[4]~q ),
	.M_bht_ptr_unfiltered_5(\M_bht_ptr_unfiltered[5]~q ),
	.M_bht_ptr_unfiltered_6(\M_bht_ptr_unfiltered[6]~q ),
	.M_bht_ptr_unfiltered_7(\M_bht_ptr_unfiltered[7]~q ),
	.F_bht_ptr_nxt_0(\F_bht_ptr_nxt[0]~combout ),
	.F_bht_ptr_nxt_1(\F_bht_ptr_nxt[1]~combout ),
	.F_bht_ptr_nxt_2(\F_bht_ptr_nxt[2]~combout ),
	.F_bht_ptr_nxt_3(\F_bht_ptr_nxt[3]~combout ),
	.F_bht_ptr_nxt_4(\F_bht_ptr_nxt[4]~combout ),
	.F_bht_ptr_nxt_5(\F_bht_ptr_nxt[5]~combout ),
	.F_bht_ptr_nxt_6(\F_bht_ptr_nxt[6]~combout ),
	.F_bht_ptr_nxt_7(\F_bht_ptr_nxt[7]~combout ),
	.M_br_mispredict(\M_br_mispredict~_wirecell_combout ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_ic_tag_module embedded_system_nios2_qsys_0_ic_tag(
	.q_b_0(\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_1(\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_7(\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_9(\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_6(\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[6] ),
	.q_b_8(\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[8] ),
	.ic_fill_valid_bits_5(\ic_fill_valid_bits[5]~q ),
	.ic_fill_valid_bits_7(\ic_fill_valid_bits[7]~q ),
	.ic_fill_valid_bits_4(\ic_fill_valid_bits[4]~q ),
	.q_b_3(\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_5(\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_2(\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_4(\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[4] ),
	.ic_fill_valid_bits_6(\ic_fill_valid_bits[6]~q ),
	.ic_fill_valid_bits_1(\ic_fill_valid_bits[1]~q ),
	.ic_fill_valid_bits_3(\ic_fill_valid_bits[3]~q ),
	.ic_fill_valid_bits_0(\ic_fill_valid_bits[0]~q ),
	.ic_fill_valid_bits_2(\ic_fill_valid_bits[2]~q ),
	.ic_fill_tag_1(ic_fill_tag_1),
	.ic_fill_tag_0(ic_fill_tag_0),
	.F_stall(\F_stall~combout ),
	.F_ic_tag_rd_addr_nxt_0(\F_ic_tag_rd_addr_nxt[0]~1_combout ),
	.F_ic_tag_rd_addr_nxt_1(\F_ic_tag_rd_addr_nxt[1]~3_combout ),
	.F_ic_tag_rd_addr_nxt_2(\F_ic_tag_rd_addr_nxt[2]~5_combout ),
	.F_ic_tag_rd_addr_nxt_3(\F_ic_tag_rd_addr_nxt[3]~7_combout ),
	.F_ic_tag_rd_addr_nxt_4(\F_ic_tag_rd_addr_nxt[4]~9_combout ),
	.F_ic_tag_rd_addr_nxt_5(\F_ic_tag_rd_addr_nxt[5]~11_combout ),
	.F_ic_tag_rd_addr_nxt_6(\F_ic_tag_rd_addr_nxt[6]~13_combout ),
	.ic_tag_wren(\ic_tag_wren~combout ),
	.ic_tag_wraddress_0(\ic_tag_wraddress[0]~q ),
	.ic_tag_wraddress_1(\ic_tag_wraddress[1]~q ),
	.ic_tag_wraddress_2(\ic_tag_wraddress[2]~q ),
	.ic_tag_wraddress_3(\ic_tag_wraddress[3]~q ),
	.ic_tag_wraddress_4(\ic_tag_wraddress[4]~q ),
	.ic_tag_wraddress_5(\ic_tag_wraddress[5]~q ),
	.ic_tag_wraddress_6(\ic_tag_wraddress[6]~q ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_ic_data_module embedded_system_nios2_qsys_0_ic_data(
	.q_b_5(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.q_b_3(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.q_b_1(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.q_b_4(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.q_b_2(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.q_b_28(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.q_b_31(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.q_b_27(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.q_b_29(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.q_b_30(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.q_b_0(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.q_b_23(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.q_b_26(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.q_b_22(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.q_b_24(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.q_b_25(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.q_b_16(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.q_b_15(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.q_b_13(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.q_b_14(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.q_b_12(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.q_b_11(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.q_b_8(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.q_b_19(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[19] ),
	.q_b_18(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[18] ),
	.q_b_17(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.q_b_10(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.q_b_9(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.q_b_21(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[21] ),
	.q_b_20(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[20] ),
	.q_b_7(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[7] ),
	.q_b_6(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[6] ),
	.ic_fill_line_6(ic_fill_line_6),
	.ic_fill_line_5(ic_fill_line_5),
	.ic_fill_line_1(ic_fill_line_1),
	.ic_fill_line_0(ic_fill_line_0),
	.ic_fill_line_4(ic_fill_line_4),
	.ic_fill_line_3(ic_fill_line_3),
	.ic_fill_line_2(ic_fill_line_2),
	.F_stall(\F_stall~combout ),
	.ic_fill_dp_offset_0(\ic_fill_dp_offset[0]~q ),
	.ic_fill_dp_offset_1(\ic_fill_dp_offset[1]~q ),
	.ic_fill_dp_offset_2(\ic_fill_dp_offset[2]~q ),
	.i_readdatavalid_d1(\i_readdatavalid_d1~q ),
	.i_readdata_d1_5(\i_readdata_d1[5]~q ),
	.F_ic_data_rd_addr_nxt_0(\F_ic_data_rd_addr_nxt[0]~3_combout ),
	.F_ic_data_rd_addr_nxt_1(\F_ic_data_rd_addr_nxt[1]~5_combout ),
	.F_ic_data_rd_addr_nxt_2(\F_ic_data_rd_addr_nxt[2]~7_combout ),
	.F_ic_tag_rd_addr_nxt_0(\F_ic_tag_rd_addr_nxt[0]~1_combout ),
	.F_ic_tag_rd_addr_nxt_1(\F_ic_tag_rd_addr_nxt[1]~3_combout ),
	.F_ic_tag_rd_addr_nxt_2(\F_ic_tag_rd_addr_nxt[2]~5_combout ),
	.F_ic_tag_rd_addr_nxt_3(\F_ic_tag_rd_addr_nxt[3]~7_combout ),
	.F_ic_tag_rd_addr_nxt_4(\F_ic_tag_rd_addr_nxt[4]~9_combout ),
	.F_ic_tag_rd_addr_nxt_5(\F_ic_tag_rd_addr_nxt[5]~11_combout ),
	.F_ic_tag_rd_addr_nxt_6(\F_ic_tag_rd_addr_nxt[6]~13_combout ),
	.i_readdata_d1_3(\i_readdata_d1[3]~q ),
	.i_readdata_d1_1(\i_readdata_d1[1]~q ),
	.i_readdata_d1_4(\i_readdata_d1[4]~q ),
	.i_readdata_d1_2(\i_readdata_d1[2]~q ),
	.i_readdata_d1_28(\i_readdata_d1[28]~q ),
	.i_readdata_d1_31(\i_readdata_d1[31]~q ),
	.i_readdata_d1_27(\i_readdata_d1[27]~q ),
	.i_readdata_d1_29(\i_readdata_d1[29]~q ),
	.i_readdata_d1_30(\i_readdata_d1[30]~q ),
	.i_readdata_d1_0(\i_readdata_d1[0]~q ),
	.i_readdata_d1_23(\i_readdata_d1[23]~q ),
	.i_readdata_d1_26(\i_readdata_d1[26]~q ),
	.i_readdata_d1_22(\i_readdata_d1[22]~q ),
	.i_readdata_d1_24(\i_readdata_d1[24]~q ),
	.i_readdata_d1_25(\i_readdata_d1[25]~q ),
	.i_readdata_d1_16(\i_readdata_d1[16]~q ),
	.i_readdata_d1_15(\i_readdata_d1[15]~q ),
	.i_readdata_d1_13(\i_readdata_d1[13]~q ),
	.i_readdata_d1_14(\i_readdata_d1[14]~q ),
	.i_readdata_d1_12(\i_readdata_d1[12]~q ),
	.i_readdata_d1_11(\i_readdata_d1[11]~q ),
	.i_readdata_d1_8(\i_readdata_d1[8]~q ),
	.i_readdata_d1_19(\i_readdata_d1[19]~q ),
	.i_readdata_d1_18(\i_readdata_d1[18]~q ),
	.i_readdata_d1_17(\i_readdata_d1[17]~q ),
	.i_readdata_d1_10(\i_readdata_d1[10]~q ),
	.i_readdata_d1_9(\i_readdata_d1[9]~q ),
	.i_readdata_d1_21(\i_readdata_d1[21]~q ),
	.i_readdata_d1_20(\i_readdata_d1[20]~q ),
	.i_readdata_d1_7(\i_readdata_d1[7]~q ),
	.i_readdata_d1_6(\i_readdata_d1[6]~q ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_nios2_oci the_embedded_system_nios2_qsys_0_nios2_oci(
	.readdata_2(readdata_2),
	.readdata_10(readdata_10),
	.readdata_18(readdata_18),
	.readdata_26(readdata_26),
	.readdata_7(readdata_7),
	.readdata_23(readdata_23),
	.readdata_15(readdata_15),
	.readdata_31(readdata_31),
	.readdata_29(readdata_29),
	.readdata_13(readdata_13),
	.readdata_28(readdata_28),
	.readdata_12(readdata_12),
	.readdata_27(readdata_27),
	.readdata_11(readdata_11),
	.readdata_25(readdata_25),
	.readdata_9(readdata_9),
	.readdata_24(readdata_24),
	.readdata_8(readdata_8),
	.readdata_6(readdata_6),
	.readdata_14(readdata_14),
	.readdata_22(readdata_22),
	.readdata_30(readdata_30),
	.readdata_5(readdata_5),
	.readdata_21(readdata_21),
	.readdata_4(readdata_4),
	.readdata_20(readdata_20),
	.readdata_3(readdata_3),
	.readdata_19(readdata_19),
	.readdata_1(readdata_1),
	.readdata_17(readdata_17),
	.readdata_0(readdata_0),
	.readdata_16(readdata_16),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.d_write(d_write),
	.saved_grant_0(saved_grant_0),
	.waitrequest(jtag_debug_module_waitrequest),
	.mem_used_1(mem_used_1),
	.hq3myc14108phmpo7y7qmhbp98hy0vq(\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.hbreak_enabled(hbreak_enabled1),
	.jtag_break(\the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_oci_debug|jtag_break~q ),
	.src0_valid(src0_valid1),
	.src1_valid(src1_valid),
	.saved_grant_1(saved_grant_1),
	.rf_source_valid(rf_source_valid),
	.r_early_rst(r_early_rst),
	.oci_single_step_mode(\the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_single_step_mode~q ),
	.address_nxt({src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.writedata_nxt({src_payload17,src_payload16,src_payload15,src_payload14,src_payload13,src_payload12,src_payload10,src_payload5,src_payload23,src_payload32,src_payload18,src_payload7,src_payload8,src_payload19,src_payload20,src_payload9,src_payload24,src_payload31,src_payload25,src_payload26,
src_payload27,src_payload21,src_payload28,src_payload29,src_payload22,src_payload30,src_payload11,src_payload6,src_payload3,src_payload4,src_payload2,src_payload}),
	.debugaccess_nxt(src_payload1),
	.byteenable_nxt({src_data_35,src_data_34,src_data_33,src_data_32}),
	.resetrequest(jtag_debug_module_resetrequest),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_1(state_1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.clk_clk(clk_clk));

dffeas \A_dc_xfer_wr_data[11] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[11]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[11]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[11] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[11] .power_up = "low";

dffeas \A_dc_xfer_wr_data[10] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[10]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[10]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[10] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[10] .power_up = "low";

dffeas \A_dc_xfer_wr_data[9] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[9]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[9]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[9] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[9] .power_up = "low";

dffeas \A_dc_xfer_wr_data[8] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[8]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[8]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[8] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[8] .power_up = "low";

dffeas \A_dc_xfer_wr_data[13] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[13]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[13]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[13] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[13] .power_up = "low";

dffeas \A_dc_xfer_wr_data[12] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[12]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[12]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[12] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[12] .power_up = "low";

dffeas \A_dc_xfer_wr_data[21] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[21]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[21]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[21] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[21] .power_up = "low";

dffeas \A_dc_xfer_wr_data[20] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[20]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[20]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[20] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[20] .power_up = "low";

dffeas \A_dc_xfer_wr_data[25] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[25]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[25]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[25] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[25] .power_up = "low";

dffeas \A_dc_xfer_wr_data[17] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[17]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[17]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[17] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[17] .power_up = "low";

dffeas \A_dc_xfer_wr_data[24] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[24]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[24]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[24] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[24] .power_up = "low";

dffeas \A_dc_xfer_wr_data[16] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[16]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[16]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[16] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[16] .power_up = "low";

dffeas \A_dc_xfer_wr_data[27] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[27]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[27]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[27] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[27] .power_up = "low";

dffeas \A_dc_xfer_wr_data[19] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[19]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[19]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[19] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[19] .power_up = "low";

dffeas \A_dc_xfer_wr_data[26] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[26]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[26]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[26] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[26] .power_up = "low";

dffeas \A_dc_xfer_wr_data[18] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[18]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[18]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[18] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[18] .power_up = "low";

dffeas \A_dc_xfer_wr_data[23] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[23]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[23]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[23] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[23] .power_up = "low";

dffeas \A_dc_xfer_wr_data[15] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[15]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[15]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[15] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[15] .power_up = "low";

dffeas \A_dc_xfer_wr_data[22] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[22]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[22]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[22] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[22] .power_up = "low";

dffeas \A_dc_xfer_wr_data[14] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[14]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[14]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[14] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[14] .power_up = "low";

dffeas \A_dc_xfer_wr_data[2] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[2]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[2]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[2] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[2] .power_up = "low";

dffeas \A_dc_xfer_wr_data[0] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[0]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[0]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[0] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[0] .power_up = "low";

dffeas \A_dc_xfer_wr_data[3] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[3]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[3]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[3] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[3] .power_up = "low";

dffeas \A_dc_xfer_wr_data[1] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[1]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[1]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[1] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[1] .power_up = "low";

dffeas \A_dc_xfer_wr_data[6] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[6]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[6]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[6] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[6] .power_up = "low";

dffeas \A_dc_xfer_wr_data[4] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[4]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[4]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[4] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[4] .power_up = "low";

dffeas \A_dc_xfer_wr_data[7] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[7]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[7]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[7] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[7] .power_up = "low";

dffeas \A_dc_xfer_wr_data[5] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[5]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[5]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[5] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[5] .power_up = "low";

dffeas \ic_fill_valid_bits[5] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[5]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[5] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[5] .power_up = "low";

dffeas \ic_fill_valid_bits[7] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[7]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[7] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[7] .power_up = "low";

dffeas \ic_fill_valid_bits[4] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[4]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[4] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[4] .power_up = "low";

dffeas \ic_fill_valid_bits[6] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[6]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[6] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[6] .power_up = "low";

dffeas \ic_fill_valid_bits[1] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[1]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[1] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[1] .power_up = "low";

dffeas \ic_fill_valid_bits[3] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[3]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[3] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[3] .power_up = "low";

dffeas \ic_fill_valid_bits[0] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[0]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[0] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[0] .power_up = "low";

dffeas \ic_fill_valid_bits[2] (
	.clk(clk_clk),
	.d(\ic_fill_valid_bits_nxt~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\ic_tag_clr_valid_bits_nxt~combout ),
	.sload(gnd),
	.ena(\ic_fill_valid_bits_en~combout ),
	.q(\ic_fill_valid_bits[2]~q ),
	.prn(vcc));
defparam \ic_fill_valid_bits[2] .is_wysiwyg = "true";
defparam \ic_fill_valid_bits[2] .power_up = "low";

dffeas \A_mul_src2[0] (
	.clk(clk_clk),
	.d(\M_src2[0]~q ),
	.asdata(\A_mul_src2[16]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[0]~q ),
	.prn(vcc));
defparam \A_mul_src2[0] .is_wysiwyg = "true";
defparam \A_mul_src2[0] .power_up = "low";

dffeas \A_mul_src2[1] (
	.clk(clk_clk),
	.d(\M_src2[1]~q ),
	.asdata(\A_mul_src2[17]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[1]~q ),
	.prn(vcc));
defparam \A_mul_src2[1] .is_wysiwyg = "true";
defparam \A_mul_src2[1] .power_up = "low";

dffeas \A_mul_src2[2] (
	.clk(clk_clk),
	.d(\M_src2[2]~q ),
	.asdata(\A_mul_src2[18]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[2]~q ),
	.prn(vcc));
defparam \A_mul_src2[2] .is_wysiwyg = "true";
defparam \A_mul_src2[2] .power_up = "low";

dffeas \A_mul_src2[3] (
	.clk(clk_clk),
	.d(\M_src2[3]~q ),
	.asdata(\A_mul_src2[19]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[3]~q ),
	.prn(vcc));
defparam \A_mul_src2[3] .is_wysiwyg = "true";
defparam \A_mul_src2[3] .power_up = "low";

dffeas \A_mul_src2[4] (
	.clk(clk_clk),
	.d(\M_src2[4]~q ),
	.asdata(\A_mul_src2[20]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[4]~q ),
	.prn(vcc));
defparam \A_mul_src2[4] .is_wysiwyg = "true";
defparam \A_mul_src2[4] .power_up = "low";

dffeas \A_mul_src2[5] (
	.clk(clk_clk),
	.d(\M_src2[5]~q ),
	.asdata(\A_mul_src2[21]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[5]~q ),
	.prn(vcc));
defparam \A_mul_src2[5] .is_wysiwyg = "true";
defparam \A_mul_src2[5] .power_up = "low";

dffeas \A_mul_src2[6] (
	.clk(clk_clk),
	.d(\M_src2[6]~q ),
	.asdata(\A_mul_src2[22]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[6]~q ),
	.prn(vcc));
defparam \A_mul_src2[6] .is_wysiwyg = "true";
defparam \A_mul_src2[6] .power_up = "low";

dffeas \A_mul_src2[7] (
	.clk(clk_clk),
	.d(\M_src2[7]~q ),
	.asdata(\A_mul_src2[23]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[7]~q ),
	.prn(vcc));
defparam \A_mul_src2[7] .is_wysiwyg = "true";
defparam \A_mul_src2[7] .power_up = "low";

dffeas \A_mul_src2[8] (
	.clk(clk_clk),
	.d(\M_src2[8]~q ),
	.asdata(\A_mul_src2[24]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[8]~q ),
	.prn(vcc));
defparam \A_mul_src2[8] .is_wysiwyg = "true";
defparam \A_mul_src2[8] .power_up = "low";

dffeas \A_mul_src2[9] (
	.clk(clk_clk),
	.d(\M_src2[9]~q ),
	.asdata(\A_mul_src2[25]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[9]~q ),
	.prn(vcc));
defparam \A_mul_src2[9] .is_wysiwyg = "true";
defparam \A_mul_src2[9] .power_up = "low";

dffeas \A_mul_src2[10] (
	.clk(clk_clk),
	.d(\M_src2[10]~q ),
	.asdata(\A_mul_src2[26]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[10]~q ),
	.prn(vcc));
defparam \A_mul_src2[10] .is_wysiwyg = "true";
defparam \A_mul_src2[10] .power_up = "low";

dffeas \A_mul_src2[11] (
	.clk(clk_clk),
	.d(\M_src2[11]~q ),
	.asdata(\A_mul_src2[27]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[11]~q ),
	.prn(vcc));
defparam \A_mul_src2[11] .is_wysiwyg = "true";
defparam \A_mul_src2[11] .power_up = "low";

dffeas \A_mul_src2[12] (
	.clk(clk_clk),
	.d(\M_src2[12]~q ),
	.asdata(\A_mul_src2[28]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[12]~q ),
	.prn(vcc));
defparam \A_mul_src2[12] .is_wysiwyg = "true";
defparam \A_mul_src2[12] .power_up = "low";

dffeas \A_mul_src2[13] (
	.clk(clk_clk),
	.d(\M_src2[13]~q ),
	.asdata(\A_mul_src2[29]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[13]~q ),
	.prn(vcc));
defparam \A_mul_src2[13] .is_wysiwyg = "true";
defparam \A_mul_src2[13] .power_up = "low";

dffeas \A_mul_src2[14] (
	.clk(clk_clk),
	.d(\M_src2[14]~q ),
	.asdata(\A_mul_src2[30]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[14]~q ),
	.prn(vcc));
defparam \A_mul_src2[14] .is_wysiwyg = "true";
defparam \A_mul_src2[14] .power_up = "low";

dffeas \A_mul_src2[15] (
	.clk(clk_clk),
	.d(\M_src2[15]~q ),
	.asdata(\A_mul_src2[31]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src2[15]~q ),
	.prn(vcc));
defparam \A_mul_src2[15] .is_wysiwyg = "true";
defparam \A_mul_src2[15] .power_up = "low";

dffeas \A_mul_src1[0] (
	.clk(clk_clk),
	.d(\M_src1[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[0]~q ),
	.prn(vcc));
defparam \A_mul_src1[0] .is_wysiwyg = "true";
defparam \A_mul_src1[0] .power_up = "low";

dffeas \A_mul_src1[1] (
	.clk(clk_clk),
	.d(\M_src1[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[1]~q ),
	.prn(vcc));
defparam \A_mul_src1[1] .is_wysiwyg = "true";
defparam \A_mul_src1[1] .power_up = "low";

dffeas \A_mul_src1[2] (
	.clk(clk_clk),
	.d(\M_src1[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[2]~q ),
	.prn(vcc));
defparam \A_mul_src1[2] .is_wysiwyg = "true";
defparam \A_mul_src1[2] .power_up = "low";

dffeas \A_mul_src1[3] (
	.clk(clk_clk),
	.d(\M_src1[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[3]~q ),
	.prn(vcc));
defparam \A_mul_src1[3] .is_wysiwyg = "true";
defparam \A_mul_src1[3] .power_up = "low";

dffeas \A_mul_src1[4] (
	.clk(clk_clk),
	.d(\M_src1[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[4]~q ),
	.prn(vcc));
defparam \A_mul_src1[4] .is_wysiwyg = "true";
defparam \A_mul_src1[4] .power_up = "low";

dffeas \A_mul_src1[5] (
	.clk(clk_clk),
	.d(\M_src1[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[5]~q ),
	.prn(vcc));
defparam \A_mul_src1[5] .is_wysiwyg = "true";
defparam \A_mul_src1[5] .power_up = "low";

dffeas \A_mul_src1[6] (
	.clk(clk_clk),
	.d(\M_src1[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[6]~q ),
	.prn(vcc));
defparam \A_mul_src1[6] .is_wysiwyg = "true";
defparam \A_mul_src1[6] .power_up = "low";

dffeas \A_mul_src1[7] (
	.clk(clk_clk),
	.d(\M_src1[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[7]~q ),
	.prn(vcc));
defparam \A_mul_src1[7] .is_wysiwyg = "true";
defparam \A_mul_src1[7] .power_up = "low";

dffeas \A_mul_src1[8] (
	.clk(clk_clk),
	.d(\M_src1[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[8]~q ),
	.prn(vcc));
defparam \A_mul_src1[8] .is_wysiwyg = "true";
defparam \A_mul_src1[8] .power_up = "low";

dffeas \A_mul_src1[9] (
	.clk(clk_clk),
	.d(\M_src1[9]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[9]~q ),
	.prn(vcc));
defparam \A_mul_src1[9] .is_wysiwyg = "true";
defparam \A_mul_src1[9] .power_up = "low";

dffeas \A_mul_src1[10] (
	.clk(clk_clk),
	.d(\M_src1[10]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[10]~q ),
	.prn(vcc));
defparam \A_mul_src1[10] .is_wysiwyg = "true";
defparam \A_mul_src1[10] .power_up = "low";

dffeas \A_mul_src1[11] (
	.clk(clk_clk),
	.d(\M_src1[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[11]~q ),
	.prn(vcc));
defparam \A_mul_src1[11] .is_wysiwyg = "true";
defparam \A_mul_src1[11] .power_up = "low";

dffeas \A_mul_src1[12] (
	.clk(clk_clk),
	.d(\M_src1[12]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[12]~q ),
	.prn(vcc));
defparam \A_mul_src1[12] .is_wysiwyg = "true";
defparam \A_mul_src1[12] .power_up = "low";

dffeas \A_mul_src1[13] (
	.clk(clk_clk),
	.d(\M_src1[13]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[13]~q ),
	.prn(vcc));
defparam \A_mul_src1[13] .is_wysiwyg = "true";
defparam \A_mul_src1[13] .power_up = "low";

dffeas \A_mul_src1[14] (
	.clk(clk_clk),
	.d(\M_src1[14]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[14]~q ),
	.prn(vcc));
defparam \A_mul_src1[14] .is_wysiwyg = "true";
defparam \A_mul_src1[14] .power_up = "low";

dffeas \A_mul_src1[15] (
	.clk(clk_clk),
	.d(\M_src1[15]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src1[15]~q ),
	.prn(vcc));
defparam \A_mul_src1[15] .is_wysiwyg = "true";
defparam \A_mul_src1[15] .power_up = "low";

dffeas \A_mul_src2[16] (
	.clk(clk_clk),
	.d(\M_src2[16]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[16]~q ),
	.prn(vcc));
defparam \A_mul_src2[16] .is_wysiwyg = "true";
defparam \A_mul_src2[16] .power_up = "low";

dffeas \A_mul_src2[17] (
	.clk(clk_clk),
	.d(\M_src2[17]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[17]~q ),
	.prn(vcc));
defparam \A_mul_src2[17] .is_wysiwyg = "true";
defparam \A_mul_src2[17] .power_up = "low";

dffeas \A_mul_src2[18] (
	.clk(clk_clk),
	.d(\M_src2[18]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[18]~q ),
	.prn(vcc));
defparam \A_mul_src2[18] .is_wysiwyg = "true";
defparam \A_mul_src2[18] .power_up = "low";

dffeas \A_mul_src2[19] (
	.clk(clk_clk),
	.d(\M_src2[19]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[19]~q ),
	.prn(vcc));
defparam \A_mul_src2[19] .is_wysiwyg = "true";
defparam \A_mul_src2[19] .power_up = "low";

dffeas \A_mul_src2[20] (
	.clk(clk_clk),
	.d(\M_src2[20]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[20]~q ),
	.prn(vcc));
defparam \A_mul_src2[20] .is_wysiwyg = "true";
defparam \A_mul_src2[20] .power_up = "low";

dffeas \A_mul_src2[21] (
	.clk(clk_clk),
	.d(\M_src2[21]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[21]~q ),
	.prn(vcc));
defparam \A_mul_src2[21] .is_wysiwyg = "true";
defparam \A_mul_src2[21] .power_up = "low";

dffeas \A_mul_src2[22] (
	.clk(clk_clk),
	.d(\M_src2[22]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[22]~q ),
	.prn(vcc));
defparam \A_mul_src2[22] .is_wysiwyg = "true";
defparam \A_mul_src2[22] .power_up = "low";

dffeas \A_mul_src2[23] (
	.clk(clk_clk),
	.d(\M_src2[23]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[23]~q ),
	.prn(vcc));
defparam \A_mul_src2[23] .is_wysiwyg = "true";
defparam \A_mul_src2[23] .power_up = "low";

dffeas \A_mul_src2[24] (
	.clk(clk_clk),
	.d(\M_src2[24]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[24]~q ),
	.prn(vcc));
defparam \A_mul_src2[24] .is_wysiwyg = "true";
defparam \A_mul_src2[24] .power_up = "low";

dffeas \A_mul_src2[25] (
	.clk(clk_clk),
	.d(\M_src2[25]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[25]~q ),
	.prn(vcc));
defparam \A_mul_src2[25] .is_wysiwyg = "true";
defparam \A_mul_src2[25] .power_up = "low";

dffeas \A_mul_src2[26] (
	.clk(clk_clk),
	.d(\M_src2[26]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[26]~q ),
	.prn(vcc));
defparam \A_mul_src2[26] .is_wysiwyg = "true";
defparam \A_mul_src2[26] .power_up = "low";

dffeas \A_mul_src2[27] (
	.clk(clk_clk),
	.d(\M_src2[27]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[27]~q ),
	.prn(vcc));
defparam \A_mul_src2[27] .is_wysiwyg = "true";
defparam \A_mul_src2[27] .power_up = "low";

dffeas \A_mul_src2[28] (
	.clk(clk_clk),
	.d(\M_src2[28]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[28]~q ),
	.prn(vcc));
defparam \A_mul_src2[28] .is_wysiwyg = "true";
defparam \A_mul_src2[28] .power_up = "low";

dffeas \A_mul_src2[29] (
	.clk(clk_clk),
	.d(\M_src2[29]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[29]~q ),
	.prn(vcc));
defparam \A_mul_src2[29] .is_wysiwyg = "true";
defparam \A_mul_src2[29] .power_up = "low";

dffeas \A_mul_src2[30] (
	.clk(clk_clk),
	.d(\M_src2[30]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[30]~q ),
	.prn(vcc));
defparam \A_mul_src2[30] .is_wysiwyg = "true";
defparam \A_mul_src2[30] .power_up = "low";

dffeas \A_mul_src2[31] (
	.clk(clk_clk),
	.d(\M_src2[31]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_mul_stall~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_src2[31]~q ),
	.prn(vcc));
defparam \A_mul_src2[31] .is_wysiwyg = "true";
defparam \A_mul_src2[31] .power_up = "low";

dffeas \A_dc_xfer_wr_data[31] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[31]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[31]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[31] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[31] .power_up = "low";

dffeas \A_dc_xfer_wr_data[29] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[29]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[29]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[29] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[29] .power_up = "low";

dffeas \A_dc_xfer_wr_data[28] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[28]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[28]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[28] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[28] .power_up = "low";

dffeas \A_dc_xfer_wr_data[30] (
	.clk(clk_clk),
	.d(\A_dc_rd_data[30]~q ),
	.asdata(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_dc_xfer_rd_data_offset_match~q ),
	.ena(vcc),
	.q(\A_dc_xfer_wr_data[30]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_data[30] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_data[30] .power_up = "low";

dffeas \A_mul_src1[16] (
	.clk(clk_clk),
	.d(\M_src1[16]~q ),
	.asdata(\A_mul_src1[0]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[16]~q ),
	.prn(vcc));
defparam \A_mul_src1[16] .is_wysiwyg = "true";
defparam \A_mul_src1[16] .power_up = "low";

dffeas \A_mul_src1[17] (
	.clk(clk_clk),
	.d(\M_src1[17]~q ),
	.asdata(\A_mul_src1[1]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[17]~q ),
	.prn(vcc));
defparam \A_mul_src1[17] .is_wysiwyg = "true";
defparam \A_mul_src1[17] .power_up = "low";

dffeas \A_mul_src1[18] (
	.clk(clk_clk),
	.d(\M_src1[18]~q ),
	.asdata(\A_mul_src1[2]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[18]~q ),
	.prn(vcc));
defparam \A_mul_src1[18] .is_wysiwyg = "true";
defparam \A_mul_src1[18] .power_up = "low";

dffeas \A_mul_src1[19] (
	.clk(clk_clk),
	.d(\M_src1[19]~q ),
	.asdata(\A_mul_src1[3]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[19]~q ),
	.prn(vcc));
defparam \A_mul_src1[19] .is_wysiwyg = "true";
defparam \A_mul_src1[19] .power_up = "low";

dffeas \A_mul_src1[20] (
	.clk(clk_clk),
	.d(\M_src1[20]~q ),
	.asdata(\A_mul_src1[4]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[20]~q ),
	.prn(vcc));
defparam \A_mul_src1[20] .is_wysiwyg = "true";
defparam \A_mul_src1[20] .power_up = "low";

dffeas \A_mul_src1[21] (
	.clk(clk_clk),
	.d(\M_src1[21]~q ),
	.asdata(\A_mul_src1[5]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[21]~q ),
	.prn(vcc));
defparam \A_mul_src1[21] .is_wysiwyg = "true";
defparam \A_mul_src1[21] .power_up = "low";

dffeas \A_mul_src1[22] (
	.clk(clk_clk),
	.d(\M_src1[22]~q ),
	.asdata(\A_mul_src1[6]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[22]~q ),
	.prn(vcc));
defparam \A_mul_src1[22] .is_wysiwyg = "true";
defparam \A_mul_src1[22] .power_up = "low";

dffeas \A_mul_src1[23] (
	.clk(clk_clk),
	.d(\M_src1[23]~q ),
	.asdata(\A_mul_src1[7]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[23]~q ),
	.prn(vcc));
defparam \A_mul_src1[23] .is_wysiwyg = "true";
defparam \A_mul_src1[23] .power_up = "low";

dffeas \A_mul_src1[24] (
	.clk(clk_clk),
	.d(\M_src1[24]~q ),
	.asdata(\A_mul_src1[8]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[24]~q ),
	.prn(vcc));
defparam \A_mul_src1[24] .is_wysiwyg = "true";
defparam \A_mul_src1[24] .power_up = "low";

dffeas \A_mul_src1[25] (
	.clk(clk_clk),
	.d(\M_src1[25]~q ),
	.asdata(\A_mul_src1[9]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[25]~q ),
	.prn(vcc));
defparam \A_mul_src1[25] .is_wysiwyg = "true";
defparam \A_mul_src1[25] .power_up = "low";

dffeas \A_mul_src1[26] (
	.clk(clk_clk),
	.d(\M_src1[26]~q ),
	.asdata(\A_mul_src1[10]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[26]~q ),
	.prn(vcc));
defparam \A_mul_src1[26] .is_wysiwyg = "true";
defparam \A_mul_src1[26] .power_up = "low";

dffeas \A_mul_src1[27] (
	.clk(clk_clk),
	.d(\M_src1[27]~q ),
	.asdata(\A_mul_src1[11]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[27]~q ),
	.prn(vcc));
defparam \A_mul_src1[27] .is_wysiwyg = "true";
defparam \A_mul_src1[27] .power_up = "low";

dffeas \A_mul_src1[28] (
	.clk(clk_clk),
	.d(\M_src1[28]~q ),
	.asdata(\A_mul_src1[12]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[28]~q ),
	.prn(vcc));
defparam \A_mul_src1[28] .is_wysiwyg = "true";
defparam \A_mul_src1[28] .power_up = "low";

dffeas \A_mul_src1[29] (
	.clk(clk_clk),
	.d(\M_src1[29]~q ),
	.asdata(\A_mul_src1[13]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[29]~q ),
	.prn(vcc));
defparam \A_mul_src1[29] .is_wysiwyg = "true";
defparam \A_mul_src1[29] .power_up = "low";

dffeas \A_mul_src1[30] (
	.clk(clk_clk),
	.d(\M_src1[30]~q ),
	.asdata(\A_mul_src1[14]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[30]~q ),
	.prn(vcc));
defparam \A_mul_src1[30] .is_wysiwyg = "true";
defparam \A_mul_src1[30] .power_up = "low";

dffeas \A_mul_src1[31] (
	.clk(clk_clk),
	.d(\M_src1[31]~q ),
	.asdata(\A_mul_src1[15]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\A_mul_stall~q ),
	.ena(vcc),
	.q(\A_mul_src1[31]~q ),
	.prn(vcc));
defparam \A_mul_src1[31] .is_wysiwyg = "true";
defparam \A_mul_src1[31] .power_up = "low";

dffeas A_dc_xfer_wr_active(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_data_active~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_wr_active~q ),
	.prn(vcc));
defparam A_dc_xfer_wr_active.is_wysiwyg = "true";
defparam A_dc_xfer_wr_active.power_up = "low";

cyclonev_lcell_comb \A_dc_wb_rd_en~0 (
	.dataa(!\A_dc_wb_rd_data_starting~q ),
	.datab(!\A_dc_wb_rd_addr_starting~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_rd_en~0 .extended_lut = "off";
defparam \A_dc_wb_rd_en~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_dc_wb_rd_en~0 .shared_arith = "off";

cyclonev_lcell_comb A_dc_wb_rd_en(
	.dataa(!hold_waitrequest),
	.datab(!d_write),
	.datac(!\A_dc_wb_wr_starting~combout ),
	.datad(!suppress_change_dest_id),
	.datae(!WideOr0),
	.dataf(!\A_dc_wb_rd_en~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_wb_rd_en.extended_lut = "off";
defparam A_dc_wb_rd_en.lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam A_dc_wb_rd_en.shared_arith = "off";

dffeas \A_dc_xfer_wr_offset[0] (
	.clk(clk_clk),
	.d(\A_dc_xfer_wr_offset_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_wr_offset[0]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_offset[0] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_offset[0] .power_up = "low";

dffeas \A_dc_xfer_wr_offset[1] (
	.clk(clk_clk),
	.d(\A_dc_xfer_wr_offset_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_wr_offset[1]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_offset[1] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_offset[1] .power_up = "low";

dffeas \A_dc_xfer_wr_offset[2] (
	.clk(clk_clk),
	.d(\A_dc_xfer_wr_offset_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_wr_offset[2]~q ),
	.prn(vcc));
defparam \A_dc_xfer_wr_offset[2] .is_wysiwyg = "true";
defparam \A_dc_xfer_wr_offset[2] .power_up = "low";

dffeas \A_dc_wb_rd_addr_offset[0] (
	.clk(clk_clk),
	.d(\A_dc_wb_rd_addr_offset_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wb_rd_en~combout ),
	.q(\A_dc_wb_rd_addr_offset[0]~q ),
	.prn(vcc));
defparam \A_dc_wb_rd_addr_offset[0] .is_wysiwyg = "true";
defparam \A_dc_wb_rd_addr_offset[0] .power_up = "low";

dffeas \A_dc_wb_rd_addr_offset[1] (
	.clk(clk_clk),
	.d(\A_dc_wb_rd_addr_offset_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wb_rd_en~combout ),
	.q(\A_dc_wb_rd_addr_offset[1]~q ),
	.prn(vcc));
defparam \A_dc_wb_rd_addr_offset[1] .is_wysiwyg = "true";
defparam \A_dc_wb_rd_addr_offset[1] .power_up = "low";

dffeas \A_dc_wb_rd_addr_offset[2] (
	.clk(clk_clk),
	.d(\A_dc_wb_rd_addr_offset_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wb_rd_en~combout ),
	.q(\A_dc_wb_rd_addr_offset[2]~q ),
	.prn(vcc));
defparam \A_dc_wb_rd_addr_offset[2] .is_wysiwyg = "true";
defparam \A_dc_wb_rd_addr_offset[2] .power_up = "low";

dffeas A_dc_fill_starting_d1(
	.clk(clk_clk),
	.d(\A_dc_fill_starting~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_fill_starting_d1~q ),
	.prn(vcc));
defparam A_dc_fill_starting_d1.is_wysiwyg = "true";
defparam A_dc_fill_starting_d1.power_up = "low";

dffeas A_en_d1(
	.clk(clk_clk),
	.d(\A_stall~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_en_d1~q ),
	.prn(vcc));
defparam A_en_d1.is_wysiwyg = "true";
defparam A_en_d1.power_up = "low";

dffeas A_ctrl_dc_index_inv(
	.clk(clk_clk),
	.d(\M_ctrl_dc_index_inv~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_dc_index_inv~q ),
	.prn(vcc));
defparam A_ctrl_dc_index_inv.is_wysiwyg = "true";
defparam A_ctrl_dc_index_inv.power_up = "low";

dffeas A_ctrl_dc_addr_inv(
	.clk(clk_clk),
	.d(\M_ctrl_dc_addr_inv~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_dc_addr_inv~q ),
	.prn(vcc));
defparam A_ctrl_dc_addr_inv.is_wysiwyg = "true";
defparam A_ctrl_dc_addr_inv.power_up = "low";

cyclonev_lcell_comb \dc_tag_wr_port_addr~0 (
	.dataa(!\A_valid~q ),
	.datab(!\A_dc_hit~q ),
	.datac(!\A_dc_fill_starting_d1~q ),
	.datad(!\A_en_d1~q ),
	.datae(!\A_ctrl_dc_index_inv~q ),
	.dataf(!\A_ctrl_dc_addr_inv~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr~0 .extended_lut = "off";
defparam \dc_tag_wr_port_addr~0 .lut_mask = 64'hFFFFFFFFFFFFFFFE;
defparam \dc_tag_wr_port_addr~0 .shared_arith = "off";

cyclonev_lcell_comb dc_tag_wr_port_en(
	.dataa(!\A_stall~combout ),
	.datab(!\M_dc_valid_st_cache_hit~0_combout ),
	.datac(!\dc_tag_wr_port_addr~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam dc_tag_wr_port_en.extended_lut = "off";
defparam dc_tag_wr_port_en.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam dc_tag_wr_port_en.shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[1]~0 (
	.dataa(!\A_mem_baddr[12]~q ),
	.datab(!\M_alu_result[12]~q ),
	.datac(!\dc_tag_wr_port_addr~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[1]~0 .extended_lut = "off";
defparam \dc_tag_wr_port_data[1]~0 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_data[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[0]~1 (
	.dataa(!\A_mem_baddr[5]~q ),
	.datab(!\M_alu_result[5]~q ),
	.datac(!\dc_tag_wr_port_addr~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[0]~1 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[0]~1 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[1]~2 (
	.dataa(!\A_mem_baddr[6]~q ),
	.datab(!\M_alu_result[6]~q ),
	.datac(!\dc_tag_wr_port_addr~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[1]~2 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[1]~2 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[2]~3 (
	.dataa(!\A_mem_baddr[7]~q ),
	.datab(!\M_alu_result[7]~q ),
	.datac(!\dc_tag_wr_port_addr~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[2]~3 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[2]~3 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[3]~4 (
	.dataa(!\A_mem_baddr[8]~q ),
	.datab(!\M_alu_result[8]~q ),
	.datac(!\dc_tag_wr_port_addr~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[3]~4 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[3]~4 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[4]~5 (
	.dataa(!\A_mem_baddr[9]~q ),
	.datab(!\M_alu_result[9]~q ),
	.datac(!\dc_tag_wr_port_addr~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[4]~5 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[4]~5 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[4]~5 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_addr[5]~6 (
	.dataa(!\A_mem_baddr[10]~q ),
	.datab(!\M_alu_result[10]~q ),
	.datac(!\dc_tag_wr_port_addr~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_addr[5]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_addr[5]~6 .extended_lut = "off";
defparam \dc_tag_wr_port_addr[5]~6 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_addr[5]~6 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[5]~q ),
	.datac(!\Add17~17_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[0]~0 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[0]~0 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[1]~1 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[6]~q ),
	.datac(!\Add17~21_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[1]~1 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[1]~1 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[2]~2 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[7]~q ),
	.datac(!\Add17~9_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[2]~2 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[2]~2 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[3]~3 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[8]~q ),
	.datac(!\Add17~1_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[3]~3 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[3]~3 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[4]~4 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[9]~q ),
	.datac(!\Add17~5_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[4]~4 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[4]~4 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_rd_port_addr[5]~5 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[10]~q ),
	.datac(!\Add17~13_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_rd_port_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_rd_port_addr[5]~5 .extended_lut = "off";
defparam \dc_tag_rd_port_addr[5]~5 .lut_mask = 64'h2727272727272727;
defparam \dc_tag_rd_port_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[2]~1 (
	.dataa(!\A_mem_baddr[13]~q ),
	.datab(!\M_alu_result[13]~q ),
	.datac(!\dc_tag_wr_port_addr~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[2]~1 .extended_lut = "off";
defparam \dc_tag_wr_port_data[2]~1 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_data[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[3]~2 (
	.dataa(!\A_valid~q ),
	.datab(!\A_dc_hit~q ),
	.datac(!\A_dc_fill_starting_d1~q ),
	.datad(!\A_en_d1~q ),
	.datae(!\A_ctrl_dc_index_inv~q ),
	.dataf(!\A_ctrl_dc_addr_inv~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[3]~2 .extended_lut = "off";
defparam \dc_tag_wr_port_data[3]~2 .lut_mask = 64'hFFFFFFFFFFFFFFEF;
defparam \dc_tag_wr_port_data[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \dc_tag_wr_port_data[0]~3 (
	.dataa(!\A_mem_baddr[11]~q ),
	.datab(!\M_alu_result[11]~q ),
	.datac(!\dc_tag_wr_port_addr~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[0]~3 .extended_lut = "off";
defparam \dc_tag_wr_port_data[0]~3 .lut_mask = 64'h5353535353535353;
defparam \dc_tag_wr_port_data[0]~3 .shared_arith = "off";

dffeas A_dc_xfer_rd_data_active(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_active~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_data_active~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_data_active.is_wysiwyg = "true";
defparam A_dc_xfer_rd_data_active.power_up = "low";

dffeas \A_dc_rd_data[11] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[11]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[11] .is_wysiwyg = "true";
defparam \A_dc_rd_data[11] .power_up = "low";

dffeas A_dc_xfer_rd_data_offset_match(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_offset_match~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_data_offset_match~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_data_offset_match.is_wysiwyg = "true";
defparam A_dc_xfer_rd_data_offset_match.power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_wr_offset_nxt[0]~0 (
	.dataa(!\A_dc_xfer_wr_offset[0]~q ),
	.datab(!\A_dc_xfer_wr_starting~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_wr_offset_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_wr_offset_nxt[0]~0 .extended_lut = "off";
defparam \A_dc_xfer_wr_offset_nxt[0]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_dc_xfer_wr_offset_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_xfer_wr_offset_nxt[1]~1 (
	.dataa(!\A_dc_xfer_wr_offset[0]~q ),
	.datab(!\A_dc_xfer_wr_offset[1]~q ),
	.datac(!\A_dc_xfer_wr_starting~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_wr_offset_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_wr_offset_nxt[1]~1 .extended_lut = "off";
defparam \A_dc_xfer_wr_offset_nxt[1]~1 .lut_mask = 64'hF6F6F6F6F6F6F6F6;
defparam \A_dc_xfer_wr_offset_nxt[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_xfer_wr_offset_nxt[2]~2 (
	.dataa(!\A_dc_xfer_wr_offset[0]~q ),
	.datab(!\A_dc_xfer_wr_offset[1]~q ),
	.datac(!\A_dc_xfer_wr_offset[2]~q ),
	.datad(!\A_dc_xfer_wr_starting~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_wr_offset_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_wr_offset_nxt[2]~2 .extended_lut = "off";
defparam \A_dc_xfer_wr_offset_nxt[2]~2 .lut_mask = 64'hFF96FF96FF96FF96;
defparam \A_dc_xfer_wr_offset_nxt[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_wb_rd_addr_offset_nxt[0]~0 (
	.dataa(!\A_dc_wb_rd_addr_starting~q ),
	.datab(!\A_dc_wb_rd_addr_offset[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_addr_offset_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_rd_addr_offset_nxt[0]~0 .extended_lut = "off";
defparam \A_dc_wb_rd_addr_offset_nxt[0]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_dc_wb_rd_addr_offset_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_wb_rd_addr_offset_nxt[1]~1 (
	.dataa(!\A_dc_wb_rd_addr_starting~q ),
	.datab(!\A_dc_wb_rd_addr_offset[0]~q ),
	.datac(!\A_dc_wb_rd_addr_offset[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_addr_offset_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_rd_addr_offset_nxt[1]~1 .extended_lut = "off";
defparam \A_dc_wb_rd_addr_offset_nxt[1]~1 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \A_dc_wb_rd_addr_offset_nxt[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_wb_rd_addr_offset_nxt[2]~2 (
	.dataa(!\A_dc_wb_rd_addr_starting~q ),
	.datab(!\A_dc_wb_rd_addr_offset[0]~q ),
	.datac(!\A_dc_wb_rd_addr_offset[1]~q ),
	.datad(!\A_dc_wb_rd_addr_offset[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_addr_offset_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_rd_addr_offset_nxt[2]~2 .extended_lut = "off";
defparam \A_dc_wb_rd_addr_offset_nxt[2]~2 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \A_dc_wb_rd_addr_offset_nxt[2]~2 .shared_arith = "off";

dffeas \A_dc_rd_data[10] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[10]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[10] .is_wysiwyg = "true";
defparam \A_dc_rd_data[10] .power_up = "low";

dffeas \A_dc_rd_data[9] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[9]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[9] .is_wysiwyg = "true";
defparam \A_dc_rd_data[9] .power_up = "low";

dffeas \A_dc_rd_data[8] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[8]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[8] .is_wysiwyg = "true";
defparam \A_dc_rd_data[8] .power_up = "low";

dffeas \A_dc_rd_data[13] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[13]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[13] .is_wysiwyg = "true";
defparam \A_dc_rd_data[13] .power_up = "low";

dffeas \A_dc_rd_data[12] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[12]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[12] .is_wysiwyg = "true";
defparam \A_dc_rd_data[12] .power_up = "low";

dffeas \A_dc_rd_data[21] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[21]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[21] .is_wysiwyg = "true";
defparam \A_dc_rd_data[21] .power_up = "low";

dffeas \A_dc_rd_data[20] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[20]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[20] .is_wysiwyg = "true";
defparam \A_dc_rd_data[20] .power_up = "low";

dffeas \A_dc_rd_data[25] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[25]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[25] .is_wysiwyg = "true";
defparam \A_dc_rd_data[25] .power_up = "low";

dffeas \A_dc_rd_data[17] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[17]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[17] .is_wysiwyg = "true";
defparam \A_dc_rd_data[17] .power_up = "low";

dffeas \A_dc_rd_data[24] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[24]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[24] .is_wysiwyg = "true";
defparam \A_dc_rd_data[24] .power_up = "low";

dffeas \A_dc_rd_data[16] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[16]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[16] .is_wysiwyg = "true";
defparam \A_dc_rd_data[16] .power_up = "low";

dffeas \A_dc_rd_data[27] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[27]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[27] .is_wysiwyg = "true";
defparam \A_dc_rd_data[27] .power_up = "low";

dffeas \A_dc_rd_data[19] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[19]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[19] .is_wysiwyg = "true";
defparam \A_dc_rd_data[19] .power_up = "low";

dffeas \A_dc_rd_data[26] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[26]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[26] .is_wysiwyg = "true";
defparam \A_dc_rd_data[26] .power_up = "low";

dffeas \A_dc_rd_data[18] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[18]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[18] .is_wysiwyg = "true";
defparam \A_dc_rd_data[18] .power_up = "low";

dffeas \A_dc_rd_data[23] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[23]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[23] .is_wysiwyg = "true";
defparam \A_dc_rd_data[23] .power_up = "low";

dffeas \A_dc_rd_data[15] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[15]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[15] .is_wysiwyg = "true";
defparam \A_dc_rd_data[15] .power_up = "low";

dffeas \A_dc_rd_data[22] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[22]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[22] .is_wysiwyg = "true";
defparam \A_dc_rd_data[22] .power_up = "low";

dffeas \A_dc_rd_data[14] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[14]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[14] .is_wysiwyg = "true";
defparam \A_dc_rd_data[14] .power_up = "low";

dffeas M_ctrl_dc_index_inv(
	.clk(clk_clk),
	.d(\E_ctrl_dc_index_inv~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_dc_index_inv~q ),
	.prn(vcc));
defparam M_ctrl_dc_index_inv.is_wysiwyg = "true";
defparam M_ctrl_dc_index_inv.power_up = "low";

dffeas M_ctrl_dc_addr_inv(
	.clk(clk_clk),
	.d(\E_ctrl_dc_addr_inv~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_dc_addr_inv~q ),
	.prn(vcc));
defparam M_ctrl_dc_addr_inv.is_wysiwyg = "true";
defparam M_ctrl_dc_addr_inv.power_up = "low";

dffeas A_valid_st_writes_mem(
	.clk(clk_clk),
	.d(\M_valid_st_writes_mem~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_valid_st_writes_mem~q ),
	.prn(vcc));
defparam A_valid_st_writes_mem.is_wysiwyg = "true";
defparam A_valid_st_writes_mem.power_up = "low";

cyclonev_lcell_comb \dc_tag_wr_port_data[4]~4 (
	.dataa(!\A_dc_fill_starting_d1~q ),
	.datab(!\dc_tag_wr_port_addr~0_combout ),
	.datac(!\A_valid_st_writes_mem~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_tag_wr_port_data[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_tag_wr_port_data[4]~4 .extended_lut = "off";
defparam \dc_tag_wr_port_data[4]~4 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \dc_tag_wr_port_data[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[22]~q ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[0]~0 .extended_lut = "off";
defparam \rf_b_rd_port_addr[0]~0 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_b_rd_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[1]~1 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[23]~q ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[1]~1 .extended_lut = "off";
defparam \rf_b_rd_port_addr[1]~1 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_b_rd_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[2]~2 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[24]~q ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[2]~2 .extended_lut = "off";
defparam \rf_b_rd_port_addr[2]~2 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_b_rd_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[3]~3 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[25]~q ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[3]~3 .extended_lut = "off";
defparam \rf_b_rd_port_addr[3]~3 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_b_rd_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \rf_b_rd_port_addr[4]~4 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[26]~q ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_b_rd_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_b_rd_port_addr[4]~4 .extended_lut = "off";
defparam \rf_b_rd_port_addr[4]~4 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_b_rd_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[27]~q ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[0]~0 .extended_lut = "off";
defparam \rf_a_rd_port_addr[0]~0 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_a_rd_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[1]~1 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[28]~q ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[1]~1 .extended_lut = "off";
defparam \rf_a_rd_port_addr[1]~1 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_a_rd_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[2]~2 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[29]~q ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[2]~2 .extended_lut = "off";
defparam \rf_a_rd_port_addr[2]~2 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_a_rd_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[3]~3 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[30]~q ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[3]~3 .extended_lut = "off";
defparam \rf_a_rd_port_addr[3]~3 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_a_rd_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \rf_a_rd_port_addr[4]~4 (
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(!\D_iw[31]~q ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\rf_a_rd_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \rf_a_rd_port_addr[4]~4 .extended_lut = "off";
defparam \rf_a_rd_port_addr[4]~4 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \rf_a_rd_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb A_dc_valid_st_bypass_hit_wr_en(
	.dataa(!\A_dc_valid_st_bypass_hit~q ),
	.datab(!\A_en_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_valid_st_bypass_hit_wr_en.extended_lut = "off";
defparam A_dc_valid_st_bypass_hit_wr_en.lut_mask = 64'h7777777777777777;
defparam A_dc_valid_st_bypass_hit_wr_en.shared_arith = "off";

cyclonev_lcell_comb dc_data_wr_port_en(
	.dataa(!\A_stall~combout ),
	.datab(!\A_dc_fill_active~q ),
	.datac(!\M_dc_valid_st_cache_hit~0_combout ),
	.datad(!\d_readdatavalid_d1~q ),
	.datae(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam dc_data_wr_port_en.extended_lut = "off";
defparam dc_data_wr_port_en.lut_mask = 64'h47FFFFFF47FFFFFF;
defparam dc_data_wr_port_en.shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[11]~0 (
	.dataa(!\M_st_data[11]~q ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[11]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[11]~0 .extended_lut = "off";
defparam \M_dc_st_data[11]~0 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[11]~0 .shared_arith = "off";

dffeas \A_dc_st_data[11] (
	.clk(clk_clk),
	.d(\M_dc_st_data[11]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[11]~q ),
	.prn(vcc));
defparam \A_dc_st_data[11] .is_wysiwyg = "true";
defparam \A_dc_st_data[11] .power_up = "low";

dffeas A_ctrl_st(
	.clk(clk_clk),
	.d(\M_ctrl_st~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_st~q ),
	.prn(vcc));
defparam A_ctrl_st.is_wysiwyg = "true";
defparam A_ctrl_st.power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[13]~0 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_byte_en[1]~q ),
	.datac(!\Equal264~0_combout ),
	.datad(!\A_dc_fill_wr_data~0_combout ),
	.datae(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.dataf(!\A_ctrl_st~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[13]~0 .extended_lut = "off";
defparam \dc_data_wr_port_data[13]~0 .lut_mask = 64'hB1FFFFFFFFFFFFFF;
defparam \dc_data_wr_port_data[13]~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_data[11]~1 (
	.dataa(!\M_dc_st_data[11]~0_combout ),
	.datab(!\A_dc_st_data[11]~q ),
	.datac(!\d_readdata_d1[11]~q ),
	.datad(!\A_st_data[11]~q ),
	.datae(!\dc_data_wr_port_data[13]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[11]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[11]~1 .extended_lut = "off";
defparam \dc_data_wr_port_data[11]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[11]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[0]~0 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[2]~q ),
	.datac(!\M_alu_result[2]~q ),
	.datad(!\A_dc_fill_dp_offset[0]~q ),
	.datae(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[0]~0 .extended_lut = "off";
defparam \dc_data_wr_port_addr[0]~0 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_wr_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[1]~1 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[3]~q ),
	.datac(!\M_alu_result[3]~q ),
	.datad(!\A_dc_fill_dp_offset[1]~q ),
	.datae(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[1]~1 .extended_lut = "off";
defparam \dc_data_wr_port_addr[1]~1 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_wr_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[2]~2 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[4]~q ),
	.datac(!\M_alu_result[4]~q ),
	.datad(!\A_dc_fill_dp_offset[2]~q ),
	.datae(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[2]~2 .extended_lut = "off";
defparam \dc_data_wr_port_addr[2]~2 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_wr_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[3]~3 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[5]~q ),
	.datac(!\M_alu_result[5]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[3]~3 .extended_lut = "off";
defparam \dc_data_wr_port_addr[3]~3 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[4]~4 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[6]~q ),
	.datac(!\M_alu_result[6]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[4]~4 .extended_lut = "off";
defparam \dc_data_wr_port_addr[4]~4 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[5]~5 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[7]~q ),
	.datac(!\M_alu_result[7]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[5]~5 .extended_lut = "off";
defparam \dc_data_wr_port_addr[5]~5 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[6]~6 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[8]~q ),
	.datac(!\M_alu_result[8]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[6]~6 .extended_lut = "off";
defparam \dc_data_wr_port_addr[6]~6 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[7]~7 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[9]~q ),
	.datac(!\M_alu_result[9]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[7]~7 .extended_lut = "off";
defparam \dc_data_wr_port_addr[7]~7 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_addr[8]~8 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[10]~q ),
	.datac(!\M_alu_result[10]~q ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_addr[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_addr[8]~8 .extended_lut = "off";
defparam \dc_data_wr_port_addr[8]~8 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \dc_data_wr_port_addr[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[0]~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[2]~q ),
	.datac(!\Add17~25_sumout ),
	.datad(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[0]~0 .extended_lut = "off";
defparam \dc_data_rd_port_addr[0]~0 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[1]~1 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[3]~q ),
	.datac(!\Add17~29_sumout ),
	.datad(!\A_dc_xfer_rd_addr_offset[1]~q ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[1]~1 .extended_lut = "off";
defparam \dc_data_rd_port_addr[1]~1 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[2]~2 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_alu_result[4]~q ),
	.datac(!\Add17~33_sumout ),
	.datad(!\A_dc_xfer_rd_addr_active~q ),
	.datae(!\A_dc_xfer_rd_addr_offset[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[2]~2 .extended_lut = "off";
defparam \dc_data_rd_port_addr[2]~2 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \dc_data_rd_port_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[3]~3 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[5]~q ),
	.datac(!\M_alu_result[5]~q ),
	.datad(!\Add17~17_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[3]~3 .extended_lut = "off";
defparam \dc_data_rd_port_addr[3]~3 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[4]~4 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[6]~q ),
	.datac(!\M_alu_result[6]~q ),
	.datad(!\Add17~21_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[4]~4 .extended_lut = "off";
defparam \dc_data_rd_port_addr[4]~4 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[5]~5 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[7]~q ),
	.datac(!\M_alu_result[7]~q ),
	.datad(!\Add17~9_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[5]~5 .extended_lut = "off";
defparam \dc_data_rd_port_addr[5]~5 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[6]~6 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[8]~q ),
	.datac(!\M_alu_result[8]~q ),
	.datad(!\Add17~1_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[6]~6 .extended_lut = "off";
defparam \dc_data_rd_port_addr[6]~6 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[7]~7 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[9]~q ),
	.datac(!\M_alu_result[9]~q ),
	.datad(!\Add17~5_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[7]~7 .extended_lut = "off";
defparam \dc_data_rd_port_addr[7]~7 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_rd_port_addr[8]~8 (
	.dataa(!\A_stall~combout ),
	.datab(!\A_mem_baddr[10]~q ),
	.datac(!\M_alu_result[10]~q ),
	.datad(!\Add17~13_sumout ),
	.datae(!\A_dc_xfer_rd_addr_active~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_rd_port_addr[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_rd_port_addr[8]~8 .extended_lut = "off";
defparam \dc_data_rd_port_addr[8]~8 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \dc_data_rd_port_addr[8]~8 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_offset_match~0 (
	.dataa(!\A_mem_baddr[2]~q ),
	.datab(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datac(!\A_valid_st_writes_mem~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_offset_match~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_offset_match~0 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_offset_match~0 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \A_dc_xfer_rd_addr_offset_match~0 .shared_arith = "off";

cyclonev_lcell_comb A_dc_xfer_rd_addr_offset_match(
	.dataa(!\A_mem_baddr[4]~q ),
	.datab(!\A_mem_baddr[3]~q ),
	.datac(!\A_dc_xfer_rd_addr_offset[1]~q ),
	.datad(!\A_dc_xfer_rd_addr_offset[2]~q ),
	.datae(!\A_dc_xfer_rd_addr_offset_match~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_offset_match~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_xfer_rd_addr_offset_match.extended_lut = "off";
defparam A_dc_xfer_rd_addr_offset_match.lut_mask = 64'h6996FFFF6996FFFF;
defparam A_dc_xfer_rd_addr_offset_match.shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[10]~1 (
	.dataa(!\M_st_data[10]~q ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[10]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[10]~1 .extended_lut = "off";
defparam \M_dc_st_data[10]~1 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[10]~1 .shared_arith = "off";

dffeas \A_dc_st_data[10] (
	.clk(clk_clk),
	.d(\M_dc_st_data[10]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[10]~q ),
	.prn(vcc));
defparam \A_dc_st_data[10] .is_wysiwyg = "true";
defparam \A_dc_st_data[10] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[10]~2 (
	.dataa(!\M_dc_st_data[10]~1_combout ),
	.datab(!\A_dc_st_data[10]~q ),
	.datac(!\d_readdata_d1[10]~q ),
	.datad(!\A_st_data[10]~q ),
	.datae(!\dc_data_wr_port_data[13]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[10]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[10]~2 .extended_lut = "off";
defparam \dc_data_wr_port_data[10]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[10]~2 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[9]~2 (
	.dataa(!\M_st_data[9]~q ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[9]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[9]~2 .extended_lut = "off";
defparam \M_dc_st_data[9]~2 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[9]~2 .shared_arith = "off";

dffeas \A_dc_st_data[9] (
	.clk(clk_clk),
	.d(\M_dc_st_data[9]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[9]~q ),
	.prn(vcc));
defparam \A_dc_st_data[9] .is_wysiwyg = "true";
defparam \A_dc_st_data[9] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[9]~3 (
	.dataa(!\M_dc_st_data[9]~2_combout ),
	.datab(!\A_dc_st_data[9]~q ),
	.datac(!\d_readdata_d1[9]~q ),
	.datad(!\A_st_data[9]~q ),
	.datae(!\dc_data_wr_port_data[13]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[9]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[9]~3 .extended_lut = "off";
defparam \dc_data_wr_port_data[9]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[9]~3 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[8]~3 (
	.dataa(!\M_st_data[8]~q ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[8]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[8]~3 .extended_lut = "off";
defparam \M_dc_st_data[8]~3 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[8]~3 .shared_arith = "off";

dffeas \A_dc_st_data[8] (
	.clk(clk_clk),
	.d(\M_dc_st_data[8]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[8]~q ),
	.prn(vcc));
defparam \A_dc_st_data[8] .is_wysiwyg = "true";
defparam \A_dc_st_data[8] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[8]~4 (
	.dataa(!\M_dc_st_data[8]~3_combout ),
	.datab(!\A_dc_st_data[8]~q ),
	.datac(!\d_readdata_d1[8]~q ),
	.datad(!\A_st_data[8]~q ),
	.datae(!\dc_data_wr_port_data[13]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[8]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[8]~4 .extended_lut = "off";
defparam \dc_data_wr_port_data[8]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[8]~4 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[13]~4 (
	.dataa(!\M_st_data[13]~q ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[13]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[13]~4 .extended_lut = "off";
defparam \M_dc_st_data[13]~4 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[13]~4 .shared_arith = "off";

dffeas \A_dc_st_data[13] (
	.clk(clk_clk),
	.d(\M_dc_st_data[13]~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[13]~q ),
	.prn(vcc));
defparam \A_dc_st_data[13] .is_wysiwyg = "true";
defparam \A_dc_st_data[13] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[13]~5 (
	.dataa(!\M_dc_st_data[13]~4_combout ),
	.datab(!\A_dc_st_data[13]~q ),
	.datac(!\d_readdata_d1[13]~q ),
	.datad(!\A_st_data[13]~q ),
	.datae(!\dc_data_wr_port_data[13]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[13]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[13]~5 .extended_lut = "off";
defparam \dc_data_wr_port_data[13]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[13]~5 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[12]~5 (
	.dataa(!\M_st_data[12]~q ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[12]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[12]~5 .extended_lut = "off";
defparam \M_dc_st_data[12]~5 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[12]~5 .shared_arith = "off";

dffeas \A_dc_st_data[12] (
	.clk(clk_clk),
	.d(\M_dc_st_data[12]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[12]~q ),
	.prn(vcc));
defparam \A_dc_st_data[12] .is_wysiwyg = "true";
defparam \A_dc_st_data[12] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[12]~6 (
	.dataa(!\M_dc_st_data[12]~5_combout ),
	.datab(!\A_dc_st_data[12]~q ),
	.datac(!\d_readdata_d1[12]~q ),
	.datad(!\A_st_data[12]~q ),
	.datae(!\dc_data_wr_port_data[13]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[12]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[12]~6 .extended_lut = "off";
defparam \dc_data_wr_port_data[12]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[12]~6 .shared_arith = "off";

dffeas \A_dc_rd_data[2] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[2]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[2] .is_wysiwyg = "true";
defparam \A_dc_rd_data[2] .power_up = "low";

dffeas \A_dc_rd_data[0] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[0]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[0] .is_wysiwyg = "true";
defparam \A_dc_rd_data[0] .power_up = "low";

dffeas \A_dc_rd_data[3] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[3]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[3] .is_wysiwyg = "true";
defparam \A_dc_rd_data[3] .power_up = "low";

dffeas \A_dc_rd_data[1] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[1]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[1] .is_wysiwyg = "true";
defparam \A_dc_rd_data[1] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[21]~6 (
	.dataa(!\M_st_data[21]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ),
	.datac(!\M_mem_byte_en[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[21]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[21]~6 .extended_lut = "off";
defparam \M_dc_st_data[21]~6 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[21]~6 .shared_arith = "off";

dffeas \A_dc_st_data[21] (
	.clk(clk_clk),
	.d(\M_dc_st_data[21]~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[21]~q ),
	.prn(vcc));
defparam \A_dc_st_data[21] .is_wysiwyg = "true";
defparam \A_dc_st_data[21] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[18]~7 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\Equal264~0_combout ),
	.datac(!\A_dc_fill_wr_data~0_combout ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(!\A_ctrl_st~q ),
	.dataf(!\A_mem_byte_en[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[18]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[18]~7 .extended_lut = "off";
defparam \dc_data_wr_port_data[18]~7 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \dc_data_wr_port_data[18]~7 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_data[21]~8 (
	.dataa(!\M_dc_st_data[21]~6_combout ),
	.datab(!\A_dc_st_data[21]~q ),
	.datac(!\d_readdata_d1[21]~q ),
	.datad(!\A_st_data[21]~q ),
	.datae(!\dc_data_wr_port_data[18]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[21]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[21]~8 .extended_lut = "off";
defparam \dc_data_wr_port_data[21]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[21]~8 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[20]~7 (
	.dataa(!\M_st_data[20]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ),
	.datac(!\M_mem_byte_en[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[20]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[20]~7 .extended_lut = "off";
defparam \M_dc_st_data[20]~7 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[20]~7 .shared_arith = "off";

dffeas \A_dc_st_data[20] (
	.clk(clk_clk),
	.d(\M_dc_st_data[20]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[20]~q ),
	.prn(vcc));
defparam \A_dc_st_data[20] .is_wysiwyg = "true";
defparam \A_dc_st_data[20] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[20]~9 (
	.dataa(!\M_dc_st_data[20]~7_combout ),
	.datab(!\A_dc_st_data[20]~q ),
	.datac(!\d_readdata_d1[20]~q ),
	.datad(!\A_st_data[20]~q ),
	.datae(!\dc_data_wr_port_data[18]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[20]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[20]~9 .extended_lut = "off";
defparam \dc_data_wr_port_data[20]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[20]~9 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[25]~8 (
	.dataa(!\M_st_data[25]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ),
	.datac(!\M_mem_byte_en[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[25]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[25]~8 .extended_lut = "off";
defparam \M_dc_st_data[25]~8 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[25]~8 .shared_arith = "off";

dffeas \A_dc_st_data[25] (
	.clk(clk_clk),
	.d(\M_dc_st_data[25]~8_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[25]~q ),
	.prn(vcc));
defparam \A_dc_st_data[25] .is_wysiwyg = "true";
defparam \A_dc_st_data[25] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[25]~10 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\Equal264~0_combout ),
	.datac(!\A_dc_fill_wr_data~0_combout ),
	.datad(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.datae(!\A_ctrl_st~q ),
	.dataf(!\A_mem_byte_en[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[25]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[25]~10 .extended_lut = "off";
defparam \dc_data_wr_port_data[25]~10 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \dc_data_wr_port_data[25]~10 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_data[25]~11 (
	.dataa(!\M_dc_st_data[25]~8_combout ),
	.datab(!\A_dc_st_data[25]~q ),
	.datac(!\d_readdata_d1[25]~q ),
	.datad(!\A_st_data[25]~q ),
	.datae(!\dc_data_wr_port_data[25]~10_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[25]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[25]~11 .extended_lut = "off";
defparam \dc_data_wr_port_data[25]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[25]~11 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[17]~9 (
	.dataa(!\M_st_data[17]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ),
	.datac(!\M_mem_byte_en[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[17]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[17]~9 .extended_lut = "off";
defparam \M_dc_st_data[17]~9 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[17]~9 .shared_arith = "off";

dffeas \A_dc_st_data[17] (
	.clk(clk_clk),
	.d(\M_dc_st_data[17]~9_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[17]~q ),
	.prn(vcc));
defparam \A_dc_st_data[17] .is_wysiwyg = "true";
defparam \A_dc_st_data[17] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[17]~12 (
	.dataa(!\M_dc_st_data[17]~9_combout ),
	.datab(!\A_dc_st_data[17]~q ),
	.datac(!\d_readdata_d1[17]~q ),
	.datad(!\A_st_data[17]~q ),
	.datae(!\dc_data_wr_port_data[18]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[17]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[17]~12 .extended_lut = "off";
defparam \dc_data_wr_port_data[17]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[17]~12 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[24]~10 (
	.dataa(!\M_st_data[24]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ),
	.datac(!\M_mem_byte_en[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[24]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[24]~10 .extended_lut = "off";
defparam \M_dc_st_data[24]~10 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[24]~10 .shared_arith = "off";

dffeas \A_dc_st_data[24] (
	.clk(clk_clk),
	.d(\M_dc_st_data[24]~10_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[24]~q ),
	.prn(vcc));
defparam \A_dc_st_data[24] .is_wysiwyg = "true";
defparam \A_dc_st_data[24] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[24]~13 (
	.dataa(!\M_dc_st_data[24]~10_combout ),
	.datab(!\A_dc_st_data[24]~q ),
	.datac(!\d_readdata_d1[24]~q ),
	.datad(!\A_st_data[24]~q ),
	.datae(!\dc_data_wr_port_data[25]~10_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[24]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[24]~13 .extended_lut = "off";
defparam \dc_data_wr_port_data[24]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[24]~13 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[16]~11 (
	.dataa(!\M_st_data[16]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ),
	.datac(!\M_mem_byte_en[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[16]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[16]~11 .extended_lut = "off";
defparam \M_dc_st_data[16]~11 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[16]~11 .shared_arith = "off";

dffeas \A_dc_st_data[16] (
	.clk(clk_clk),
	.d(\M_dc_st_data[16]~11_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[16]~q ),
	.prn(vcc));
defparam \A_dc_st_data[16] .is_wysiwyg = "true";
defparam \A_dc_st_data[16] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[16]~14 (
	.dataa(!\M_dc_st_data[16]~11_combout ),
	.datab(!\A_dc_st_data[16]~q ),
	.datac(!\d_readdata_d1[16]~q ),
	.datad(!\A_st_data[16]~q ),
	.datae(!\dc_data_wr_port_data[18]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[16]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[16]~14 .extended_lut = "off";
defparam \dc_data_wr_port_data[16]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[16]~14 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[27]~12 (
	.dataa(!\M_st_data[27]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ),
	.datac(!\M_mem_byte_en[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[27]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[27]~12 .extended_lut = "off";
defparam \M_dc_st_data[27]~12 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[27]~12 .shared_arith = "off";

dffeas \A_dc_st_data[27] (
	.clk(clk_clk),
	.d(\M_dc_st_data[27]~12_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[27]~q ),
	.prn(vcc));
defparam \A_dc_st_data[27] .is_wysiwyg = "true";
defparam \A_dc_st_data[27] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[27]~15 (
	.dataa(!\M_dc_st_data[27]~12_combout ),
	.datab(!\A_dc_st_data[27]~q ),
	.datac(!\d_readdata_d1[27]~q ),
	.datad(!\A_st_data[27]~q ),
	.datae(!\dc_data_wr_port_data[25]~10_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[27]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[27]~15 .extended_lut = "off";
defparam \dc_data_wr_port_data[27]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[27]~15 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[19]~13 (
	.dataa(!\M_st_data[19]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ),
	.datac(!\M_mem_byte_en[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[19]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[19]~13 .extended_lut = "off";
defparam \M_dc_st_data[19]~13 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[19]~13 .shared_arith = "off";

dffeas \A_dc_st_data[19] (
	.clk(clk_clk),
	.d(\M_dc_st_data[19]~13_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[19]~q ),
	.prn(vcc));
defparam \A_dc_st_data[19] .is_wysiwyg = "true";
defparam \A_dc_st_data[19] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[19]~16 (
	.dataa(!\M_dc_st_data[19]~13_combout ),
	.datab(!\A_dc_st_data[19]~q ),
	.datac(!\d_readdata_d1[19]~q ),
	.datad(!\A_st_data[19]~q ),
	.datae(!\dc_data_wr_port_data[18]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[19]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[19]~16 .extended_lut = "off";
defparam \dc_data_wr_port_data[19]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[19]~16 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[26]~14 (
	.dataa(!\M_st_data[26]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ),
	.datac(!\M_mem_byte_en[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[26]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[26]~14 .extended_lut = "off";
defparam \M_dc_st_data[26]~14 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[26]~14 .shared_arith = "off";

dffeas \A_dc_st_data[26] (
	.clk(clk_clk),
	.d(\M_dc_st_data[26]~14_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[26]~q ),
	.prn(vcc));
defparam \A_dc_st_data[26] .is_wysiwyg = "true";
defparam \A_dc_st_data[26] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[26]~17 (
	.dataa(!\M_dc_st_data[26]~14_combout ),
	.datab(!\A_dc_st_data[26]~q ),
	.datac(!\d_readdata_d1[26]~q ),
	.datad(!\A_st_data[26]~q ),
	.datae(!\dc_data_wr_port_data[25]~10_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[26]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[26]~17 .extended_lut = "off";
defparam \dc_data_wr_port_data[26]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[26]~17 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[18]~15 (
	.dataa(!\M_st_data[18]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ),
	.datac(!\M_mem_byte_en[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[18]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[18]~15 .extended_lut = "off";
defparam \M_dc_st_data[18]~15 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[18]~15 .shared_arith = "off";

dffeas \A_dc_st_data[18] (
	.clk(clk_clk),
	.d(\M_dc_st_data[18]~15_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[18]~q ),
	.prn(vcc));
defparam \A_dc_st_data[18] .is_wysiwyg = "true";
defparam \A_dc_st_data[18] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[18]~18 (
	.dataa(!\M_dc_st_data[18]~15_combout ),
	.datab(!\A_dc_st_data[18]~q ),
	.datac(!\d_readdata_d1[18]~q ),
	.datad(!\A_st_data[18]~q ),
	.datae(!\dc_data_wr_port_data[18]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[18]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[18]~18 .extended_lut = "off";
defparam \dc_data_wr_port_data[18]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[18]~18 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[23]~16 (
	.dataa(!\M_st_data[23]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\M_mem_byte_en[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[23]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[23]~16 .extended_lut = "off";
defparam \M_dc_st_data[23]~16 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[23]~16 .shared_arith = "off";

dffeas \A_dc_st_data[23] (
	.clk(clk_clk),
	.d(\M_dc_st_data[23]~16_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[23]~q ),
	.prn(vcc));
defparam \A_dc_st_data[23] .is_wysiwyg = "true";
defparam \A_dc_st_data[23] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[23]~19 (
	.dataa(!\M_dc_st_data[23]~16_combout ),
	.datab(!\A_dc_st_data[23]~q ),
	.datac(!\d_readdata_d1[23]~q ),
	.datad(!\A_st_data[23]~q ),
	.datae(!\dc_data_wr_port_data[18]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[23]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[23]~19 .extended_lut = "off";
defparam \dc_data_wr_port_data[23]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[23]~19 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[15]~17 (
	.dataa(!\M_st_data[15]~q ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[15]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[15]~17 .extended_lut = "off";
defparam \M_dc_st_data[15]~17 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[15]~17 .shared_arith = "off";

dffeas \A_dc_st_data[15] (
	.clk(clk_clk),
	.d(\M_dc_st_data[15]~17_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[15]~q ),
	.prn(vcc));
defparam \A_dc_st_data[15] .is_wysiwyg = "true";
defparam \A_dc_st_data[15] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[15]~20 (
	.dataa(!\M_dc_st_data[15]~17_combout ),
	.datab(!\A_dc_st_data[15]~q ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\A_st_data[15]~q ),
	.datae(!\dc_data_wr_port_data[13]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[15]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[15]~20 .extended_lut = "off";
defparam \dc_data_wr_port_data[15]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[15]~20 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[22]~18 (
	.dataa(!\M_st_data[22]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ),
	.datac(!\M_mem_byte_en[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[22]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[22]~18 .extended_lut = "off";
defparam \M_dc_st_data[22]~18 .lut_mask = 64'h5353535353535353;
defparam \M_dc_st_data[22]~18 .shared_arith = "off";

dffeas \A_dc_st_data[22] (
	.clk(clk_clk),
	.d(\M_dc_st_data[22]~18_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[22]~q ),
	.prn(vcc));
defparam \A_dc_st_data[22] .is_wysiwyg = "true";
defparam \A_dc_st_data[22] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[22]~21 (
	.dataa(!\M_dc_st_data[22]~18_combout ),
	.datab(!\A_dc_st_data[22]~q ),
	.datac(!\d_readdata_d1[22]~q ),
	.datad(!\A_st_data[22]~q ),
	.datae(!\dc_data_wr_port_data[18]~7_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[22]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[22]~21 .extended_lut = "off";
defparam \dc_data_wr_port_data[22]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[22]~21 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[14]~19 (
	.dataa(!\M_st_data[14]~q ),
	.datab(!\M_mem_byte_en[1]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[14]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[14]~19 .extended_lut = "off";
defparam \M_dc_st_data[14]~19 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[14]~19 .shared_arith = "off";

dffeas \A_dc_st_data[14] (
	.clk(clk_clk),
	.d(\M_dc_st_data[14]~19_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[14]~q ),
	.prn(vcc));
defparam \A_dc_st_data[14] .is_wysiwyg = "true";
defparam \A_dc_st_data[14] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[14]~22 (
	.dataa(!\M_dc_st_data[14]~19_combout ),
	.datab(!\A_dc_st_data[14]~q ),
	.datac(!\d_readdata_d1[14]~q ),
	.datad(!\A_st_data[14]~q ),
	.datae(!\dc_data_wr_port_data[13]~0_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[14]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[14]~22 .extended_lut = "off";
defparam \dc_data_wr_port_data[14]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[14]~22 .shared_arith = "off";

dffeas \i_readdata_d1[5] (
	.clk(clk_clk),
	.d(i_readdata[5]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[5]~q ),
	.prn(vcc));
defparam \i_readdata_d1[5] .is_wysiwyg = "true";
defparam \i_readdata_d1[5] .power_up = "low";

dffeas \i_readdata_d1[3] (
	.clk(clk_clk),
	.d(i_readdata[3]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[3]~q ),
	.prn(vcc));
defparam \i_readdata_d1[3] .is_wysiwyg = "true";
defparam \i_readdata_d1[3] .power_up = "low";

dffeas \i_readdata_d1[1] (
	.clk(clk_clk),
	.d(i_readdata[1]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[1]~q ),
	.prn(vcc));
defparam \i_readdata_d1[1] .is_wysiwyg = "true";
defparam \i_readdata_d1[1] .power_up = "low";

dffeas \i_readdata_d1[4] (
	.clk(clk_clk),
	.d(i_readdata[4]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[4]~q ),
	.prn(vcc));
defparam \i_readdata_d1[4] .is_wysiwyg = "true";
defparam \i_readdata_d1[4] .power_up = "low";

dffeas \i_readdata_d1[2] (
	.clk(clk_clk),
	.d(i_readdata[2]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[2]~q ),
	.prn(vcc));
defparam \i_readdata_d1[2] .is_wysiwyg = "true";
defparam \i_readdata_d1[2] .power_up = "low";

dffeas \i_readdata_d1[28] (
	.clk(clk_clk),
	.d(i_readdata[28]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[28]~q ),
	.prn(vcc));
defparam \i_readdata_d1[28] .is_wysiwyg = "true";
defparam \i_readdata_d1[28] .power_up = "low";

dffeas \i_readdata_d1[31] (
	.clk(clk_clk),
	.d(i_readdata[31]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[31]~q ),
	.prn(vcc));
defparam \i_readdata_d1[31] .is_wysiwyg = "true";
defparam \i_readdata_d1[31] .power_up = "low";

dffeas \i_readdata_d1[27] (
	.clk(clk_clk),
	.d(i_readdata[27]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[27]~q ),
	.prn(vcc));
defparam \i_readdata_d1[27] .is_wysiwyg = "true";
defparam \i_readdata_d1[27] .power_up = "low";

dffeas \i_readdata_d1[29] (
	.clk(clk_clk),
	.d(i_readdata[29]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[29]~q ),
	.prn(vcc));
defparam \i_readdata_d1[29] .is_wysiwyg = "true";
defparam \i_readdata_d1[29] .power_up = "low";

dffeas \i_readdata_d1[30] (
	.clk(clk_clk),
	.d(i_readdata[30]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[30]~q ),
	.prn(vcc));
defparam \i_readdata_d1[30] .is_wysiwyg = "true";
defparam \i_readdata_d1[30] .power_up = "low";

dffeas \i_readdata_d1[0] (
	.clk(clk_clk),
	.d(i_readdata[0]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[0]~q ),
	.prn(vcc));
defparam \i_readdata_d1[0] .is_wysiwyg = "true";
defparam \i_readdata_d1[0] .power_up = "low";

dffeas \i_readdata_d1[23] (
	.clk(clk_clk),
	.d(i_readdata[23]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[23]~q ),
	.prn(vcc));
defparam \i_readdata_d1[23] .is_wysiwyg = "true";
defparam \i_readdata_d1[23] .power_up = "low";

dffeas \i_readdata_d1[26] (
	.clk(clk_clk),
	.d(i_readdata[26]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[26]~q ),
	.prn(vcc));
defparam \i_readdata_d1[26] .is_wysiwyg = "true";
defparam \i_readdata_d1[26] .power_up = "low";

dffeas \i_readdata_d1[22] (
	.clk(clk_clk),
	.d(i_readdata[22]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[22]~q ),
	.prn(vcc));
defparam \i_readdata_d1[22] .is_wysiwyg = "true";
defparam \i_readdata_d1[22] .power_up = "low";

dffeas \i_readdata_d1[24] (
	.clk(clk_clk),
	.d(i_readdata[24]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[24]~q ),
	.prn(vcc));
defparam \i_readdata_d1[24] .is_wysiwyg = "true";
defparam \i_readdata_d1[24] .power_up = "low";

dffeas \i_readdata_d1[25] (
	.clk(clk_clk),
	.d(i_readdata[25]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[25]~q ),
	.prn(vcc));
defparam \i_readdata_d1[25] .is_wysiwyg = "true";
defparam \i_readdata_d1[25] .power_up = "low";

dffeas ic_tag_clr_valid_bits(
	.clk(clk_clk),
	.d(\ic_tag_clr_valid_bits~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_clr_valid_bits~q ),
	.prn(vcc));
defparam ic_tag_clr_valid_bits.is_wysiwyg = "true";
defparam ic_tag_clr_valid_bits.power_up = "low";

cyclonev_lcell_comb ic_tag_wren(
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\ic_tag_clr_valid_bits~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wren~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_tag_wren.extended_lut = "off";
defparam ic_tag_wren.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam ic_tag_wren.shared_arith = "off";

dffeas \ic_tag_wraddress[0] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[0]~8_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[0]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[0] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[0] .power_up = "low";

dffeas \ic_tag_wraddress[1] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[1]~10_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[1]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[1] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[1] .power_up = "low";

dffeas \ic_tag_wraddress[2] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[2]~11_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[2]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[2] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[2] .power_up = "low";

dffeas \ic_tag_wraddress[3] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[3]~12_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[3]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[3] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[3] .power_up = "low";

dffeas \ic_tag_wraddress[4] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[4]~13_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[4]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[4] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[4] .power_up = "low";

dffeas \ic_tag_wraddress[5] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[5]~14_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[5]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[5] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[5] .power_up = "low";

dffeas \ic_tag_wraddress[6] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt[6]~15_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_tag_wraddress[6]~q ),
	.prn(vcc));
defparam \ic_tag_wraddress[6] .is_wysiwyg = "true";
defparam \ic_tag_wraddress[6] .power_up = "low";

dffeas \i_readdata_d1[16] (
	.clk(clk_clk),
	.d(i_readdata[16]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[16]~q ),
	.prn(vcc));
defparam \i_readdata_d1[16] .is_wysiwyg = "true";
defparam \i_readdata_d1[16] .power_up = "low";

dffeas \i_readdata_d1[15] (
	.clk(clk_clk),
	.d(i_readdata[15]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[15]~q ),
	.prn(vcc));
defparam \i_readdata_d1[15] .is_wysiwyg = "true";
defparam \i_readdata_d1[15] .power_up = "low";

dffeas \i_readdata_d1[13] (
	.clk(clk_clk),
	.d(i_readdata[13]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[13]~q ),
	.prn(vcc));
defparam \i_readdata_d1[13] .is_wysiwyg = "true";
defparam \i_readdata_d1[13] .power_up = "low";

dffeas \i_readdata_d1[14] (
	.clk(clk_clk),
	.d(i_readdata[14]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[14]~q ),
	.prn(vcc));
defparam \i_readdata_d1[14] .is_wysiwyg = "true";
defparam \i_readdata_d1[14] .power_up = "low";

dffeas \i_readdata_d1[12] (
	.clk(clk_clk),
	.d(i_readdata[12]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[12]~q ),
	.prn(vcc));
defparam \i_readdata_d1[12] .is_wysiwyg = "true";
defparam \i_readdata_d1[12] .power_up = "low";

dffeas \i_readdata_d1[11] (
	.clk(clk_clk),
	.d(i_readdata[11]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[11]~q ),
	.prn(vcc));
defparam \i_readdata_d1[11] .is_wysiwyg = "true";
defparam \i_readdata_d1[11] .power_up = "low";

cyclonev_lcell_comb \E_ctrl_dc_index_inv~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[4]~q ),
	.datad(!\E_iw[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_dc_index_inv~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_dc_index_inv~0 .extended_lut = "off";
defparam \E_ctrl_dc_index_inv~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_ctrl_dc_index_inv~0 .shared_arith = "off";

dffeas M_ctrl_st(
	.clk(clk_clk),
	.d(\M_ctrl_st_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_st~q ),
	.prn(vcc));
defparam M_ctrl_st.is_wysiwyg = "true";
defparam M_ctrl_st.power_up = "low";

cyclonev_lcell_comb M_valid_st_writes_mem(
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_st~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_valid_st_writes_mem~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_valid_st_writes_mem.extended_lut = "off";
defparam M_valid_st_writes_mem.lut_mask = 64'h7777777777777777;
defparam M_valid_st_writes_mem.shared_arith = "off";

dffeas \i_readdata_d1[8] (
	.clk(clk_clk),
	.d(i_readdata[8]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[8]~q ),
	.prn(vcc));
defparam \i_readdata_d1[8] .is_wysiwyg = "true";
defparam \i_readdata_d1[8] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[2]~20 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\M_st_data[2]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[2]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[2]~20 .extended_lut = "off";
defparam \M_dc_st_data[2]~20 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[2]~20 .shared_arith = "off";

dffeas \A_dc_st_data[2] (
	.clk(clk_clk),
	.d(\M_dc_st_data[2]~20_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[2]~q ),
	.prn(vcc));
defparam \A_dc_st_data[2] .is_wysiwyg = "true";
defparam \A_dc_st_data[2] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[1]~23 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_byte_en[0]~q ),
	.datac(!\Equal264~0_combout ),
	.datad(!\A_dc_fill_wr_data~0_combout ),
	.datae(!\A_dc_valid_st_bypass_hit_wr_en~combout ),
	.dataf(!\A_ctrl_st~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[1]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[1]~23 .extended_lut = "off";
defparam \dc_data_wr_port_data[1]~23 .lut_mask = 64'hB1FFFFFFFFFFFFFF;
defparam \dc_data_wr_port_data[1]~23 .shared_arith = "off";

cyclonev_lcell_comb \dc_data_wr_port_data[2]~24 (
	.dataa(!\M_dc_st_data[2]~20_combout ),
	.datab(!\A_dc_st_data[2]~q ),
	.datac(!\d_readdata_d1[2]~q ),
	.datad(!\A_st_data[2]~q ),
	.datae(!\dc_data_wr_port_data[1]~23_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[2]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[2]~24 .extended_lut = "off";
defparam \dc_data_wr_port_data[2]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[2]~24 .shared_arith = "off";

dffeas M_ctrl_br_cond(
	.clk(clk_clk),
	.d(\E_ctrl_br_cond~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_br_cond~q ),
	.prn(vcc));
defparam M_ctrl_br_cond.is_wysiwyg = "true";
defparam M_ctrl_br_cond.power_up = "low";

cyclonev_lcell_comb M_bht_wr_en_unfiltered(
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_br_cond~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_bht_wr_en_unfiltered~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_bht_wr_en_unfiltered.extended_lut = "off";
defparam M_bht_wr_en_unfiltered.lut_mask = 64'h7777777777777777;
defparam M_bht_wr_en_unfiltered.shared_arith = "off";

dffeas \M_bht_data[1] (
	.clk(clk_clk),
	.d(\E_bht_data[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_data[1]~q ),
	.prn(vcc));
defparam \M_bht_data[1] .is_wysiwyg = "true";
defparam \M_bht_data[1] .power_up = "low";

dffeas \M_bht_data[0] (
	.clk(clk_clk),
	.d(\E_bht_data[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_data[0]~q ),
	.prn(vcc));
defparam \M_bht_data[0] .is_wysiwyg = "true";
defparam \M_bht_data[0] .power_up = "low";

dffeas M_br_mispredict(
	.clk(clk_clk),
	.d(\E_br_mispredict~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_br_mispredict~q ),
	.prn(vcc));
defparam M_br_mispredict.is_wysiwyg = "true";
defparam M_br_mispredict.power_up = "low";

cyclonev_lcell_comb \M_bht_wr_data_unfiltered[1]~0 (
	.dataa(!\M_bht_data[1]~q ),
	.datab(!\M_bht_data[0]~q ),
	.datac(!\M_br_mispredict~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_bht_wr_data_unfiltered[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_bht_wr_data_unfiltered[1]~0 .extended_lut = "off";
defparam \M_bht_wr_data_unfiltered[1]~0 .lut_mask = 64'h9696969696969696;
defparam \M_bht_wr_data_unfiltered[1]~0 .shared_arith = "off";

dffeas \M_bht_ptr_unfiltered[0] (
	.clk(clk_clk),
	.d(\E_bht_ptr[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[0]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[0] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[0] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[1] (
	.clk(clk_clk),
	.d(\E_bht_ptr[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[1]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[1] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[1] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[2] (
	.clk(clk_clk),
	.d(\E_bht_ptr[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[2]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[2] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[2] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[3] (
	.clk(clk_clk),
	.d(\E_bht_ptr[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[3]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[3] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[3] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[4] (
	.clk(clk_clk),
	.d(\E_bht_ptr[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[4]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[4] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[4] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[5] (
	.clk(clk_clk),
	.d(\E_bht_ptr[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[5]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[5] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[5] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[6] (
	.clk(clk_clk),
	.d(\E_bht_ptr[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[6]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[6] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[6] .power_up = "low";

dffeas \M_bht_ptr_unfiltered[7] (
	.clk(clk_clk),
	.d(\E_bht_ptr[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_bht_ptr_unfiltered[7]~q ),
	.prn(vcc));
defparam \M_bht_ptr_unfiltered[7] .is_wysiwyg = "true";
defparam \M_bht_ptr_unfiltered[7] .power_up = "low";

dffeas \M_br_cond_taken_history[0] (
	.clk(clk_clk),
	.d(\E_br_result~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~1_combout ),
	.q(\M_br_cond_taken_history[0]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[0] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[0] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[0] (
	.dataa(!\E_src1[2]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~2_combout ),
	.dataf(!\M_br_cond_taken_history[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[0] .extended_lut = "off";
defparam \F_bht_ptr_nxt[0] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[0] .shared_arith = "off";

dffeas \M_br_cond_taken_history[1] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~1_combout ),
	.q(\M_br_cond_taken_history[1]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[1] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[1] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[1] (
	.dataa(!\E_src1[3]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[1]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[1]~4_combout ),
	.dataf(!\M_br_cond_taken_history[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[1] .extended_lut = "off";
defparam \F_bht_ptr_nxt[1] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[1] .shared_arith = "off";

dffeas \M_br_cond_taken_history[2] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~1_combout ),
	.q(\M_br_cond_taken_history[2]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[2] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[2] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[2] (
	.dataa(!\E_src1[4]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[2]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~6_combout ),
	.dataf(!\M_br_cond_taken_history[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[2] .extended_lut = "off";
defparam \F_bht_ptr_nxt[2] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[2] .shared_arith = "off";

dffeas \M_br_cond_taken_history[3] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~1_combout ),
	.q(\M_br_cond_taken_history[3]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[3] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[3] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[3] (
	.dataa(!\E_src1[5]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[3]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[0]~0_combout ),
	.dataf(!\M_br_cond_taken_history[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[3] .extended_lut = "off";
defparam \F_bht_ptr_nxt[3] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[3] .shared_arith = "off";

dffeas \M_br_cond_taken_history[4] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~1_combout ),
	.q(\M_br_cond_taken_history[4]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[4] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[4] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[4] (
	.dataa(!\E_src1[6]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[4]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[1]~2_combout ),
	.dataf(!\M_br_cond_taken_history[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[4] .extended_lut = "off";
defparam \F_bht_ptr_nxt[4] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[4] .shared_arith = "off";

dffeas \M_br_cond_taken_history[5] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~1_combout ),
	.q(\M_br_cond_taken_history[5]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[5] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[5] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[5] (
	.dataa(!\E_src1[7]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[5]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[2]~4_combout ),
	.dataf(!\M_br_cond_taken_history[5]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[5] .extended_lut = "off";
defparam \F_bht_ptr_nxt[5] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[5] .shared_arith = "off";

dffeas \M_br_cond_taken_history[6] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~1_combout ),
	.q(\M_br_cond_taken_history[6]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[6] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[6] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[6] (
	.dataa(!\E_src1[8]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[6]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~6_combout ),
	.dataf(!\M_br_cond_taken_history[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[6] .extended_lut = "off";
defparam \F_bht_ptr_nxt[6] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[6] .shared_arith = "off";

dffeas \M_br_cond_taken_history[7] (
	.clk(clk_clk),
	.d(\M_br_cond_taken_history[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\M_br_cond_taken_history[0]~1_combout ),
	.q(\M_br_cond_taken_history[7]~q ),
	.prn(vcc));
defparam \M_br_cond_taken_history[7] .is_wysiwyg = "true";
defparam \M_br_cond_taken_history[7] .power_up = "low";

cyclonev_lcell_comb \F_bht_ptr_nxt[7] (
	.dataa(!\E_src1[9]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[7]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[4]~8_combout ),
	.dataf(!\M_br_cond_taken_history[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_bht_ptr_nxt[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_bht_ptr_nxt[7] .extended_lut = "off";
defparam \F_bht_ptr_nxt[7] .lut_mask = 64'h6996966996696996;
defparam \F_bht_ptr_nxt[7] .shared_arith = "off";

dffeas \i_readdata_d1[19] (
	.clk(clk_clk),
	.d(i_readdata[19]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[19]~q ),
	.prn(vcc));
defparam \i_readdata_d1[19] .is_wysiwyg = "true";
defparam \i_readdata_d1[19] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[29]~21 (
	.dataa(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[29]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[29]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[29]~21 .extended_lut = "off";
defparam \M_dc_st_data[29]~21 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[29]~21 .shared_arith = "off";

dffeas \A_dc_st_data[29] (
	.clk(clk_clk),
	.d(\M_dc_st_data[29]~21_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[29]~q ),
	.prn(vcc));
defparam \A_dc_st_data[29] .is_wysiwyg = "true";
defparam \A_dc_st_data[29] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[29]~25 (
	.dataa(!\M_dc_st_data[29]~21_combout ),
	.datab(!\A_dc_st_data[29]~q ),
	.datac(!\d_readdata_d1[29]~q ),
	.datad(!\A_st_data[29]~q ),
	.datae(!\dc_data_wr_port_data[25]~10_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[29]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[29]~25 .extended_lut = "off";
defparam \dc_data_wr_port_data[29]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[29]~25 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[7]~22 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\M_st_data[7]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[7]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[7]~22 .extended_lut = "off";
defparam \M_dc_st_data[7]~22 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[7]~22 .shared_arith = "off";

dffeas \A_dc_st_data[7] (
	.clk(clk_clk),
	.d(\M_dc_st_data[7]~22_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[7]~q ),
	.prn(vcc));
defparam \A_dc_st_data[7] .is_wysiwyg = "true";
defparam \A_dc_st_data[7] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[7]~26 (
	.dataa(!\M_dc_st_data[7]~22_combout ),
	.datab(!\A_dc_st_data[7]~q ),
	.datac(!\d_readdata_d1[7]~q ),
	.datad(!\A_st_data[7]~q ),
	.datae(!\dc_data_wr_port_data[1]~23_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[7]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[7]~26 .extended_lut = "off";
defparam \dc_data_wr_port_data[7]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[7]~26 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[31]~23 (
	.dataa(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[31]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[31]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[31]~23 .extended_lut = "off";
defparam \M_dc_st_data[31]~23 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[31]~23 .shared_arith = "off";

dffeas \A_dc_st_data[31] (
	.clk(clk_clk),
	.d(\M_dc_st_data[31]~23_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[31]~q ),
	.prn(vcc));
defparam \A_dc_st_data[31] .is_wysiwyg = "true";
defparam \A_dc_st_data[31] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[31]~27 (
	.dataa(!\M_dc_st_data[31]~23_combout ),
	.datab(!\A_dc_st_data[31]~q ),
	.datac(!\d_readdata_d1[31]~q ),
	.datad(!\A_st_data[31]~q ),
	.datae(!\dc_data_wr_port_data[25]~10_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[31]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[31]~27 .extended_lut = "off";
defparam \dc_data_wr_port_data[31]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[31]~27 .shared_arith = "off";

dffeas \i_readdata_d1[18] (
	.clk(clk_clk),
	.d(i_readdata[18]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[18]~q ),
	.prn(vcc));
defparam \i_readdata_d1[18] .is_wysiwyg = "true";
defparam \i_readdata_d1[18] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[28]~24 (
	.dataa(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[28]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[28]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[28]~24 .extended_lut = "off";
defparam \M_dc_st_data[28]~24 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[28]~24 .shared_arith = "off";

dffeas \A_dc_st_data[28] (
	.clk(clk_clk),
	.d(\M_dc_st_data[28]~24_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[28]~q ),
	.prn(vcc));
defparam \A_dc_st_data[28] .is_wysiwyg = "true";
defparam \A_dc_st_data[28] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[28]~28 (
	.dataa(!\M_dc_st_data[28]~24_combout ),
	.datab(!\A_dc_st_data[28]~q ),
	.datac(!\d_readdata_d1[28]~q ),
	.datad(!\A_st_data[28]~q ),
	.datae(!\dc_data_wr_port_data[25]~10_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[28]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[28]~28 .extended_lut = "off";
defparam \dc_data_wr_port_data[28]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[28]~28 .shared_arith = "off";

dffeas \i_readdata_d1[17] (
	.clk(clk_clk),
	.d(i_readdata[17]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[17]~q ),
	.prn(vcc));
defparam \i_readdata_d1[17] .is_wysiwyg = "true";
defparam \i_readdata_d1[17] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[6]~25 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\M_st_data[6]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[6]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[6]~25 .extended_lut = "off";
defparam \M_dc_st_data[6]~25 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[6]~25 .shared_arith = "off";

dffeas \A_dc_st_data[6] (
	.clk(clk_clk),
	.d(\M_dc_st_data[6]~25_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[6]~q ),
	.prn(vcc));
defparam \A_dc_st_data[6] .is_wysiwyg = "true";
defparam \A_dc_st_data[6] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[6]~29 (
	.dataa(!\M_dc_st_data[6]~25_combout ),
	.datab(!\A_dc_st_data[6]~q ),
	.datac(!\d_readdata_d1[6]~q ),
	.datad(!\A_st_data[6]~q ),
	.datae(!\dc_data_wr_port_data[1]~23_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[6]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[6]~29 .extended_lut = "off";
defparam \dc_data_wr_port_data[6]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[6]~29 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[30]~26 (
	.dataa(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ),
	.datab(!\M_mem_byte_en[3]~q ),
	.datac(!\M_st_data[30]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[30]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[30]~26 .extended_lut = "off";
defparam \M_dc_st_data[30]~26 .lut_mask = 64'h4747474747474747;
defparam \M_dc_st_data[30]~26 .shared_arith = "off";

dffeas \A_dc_st_data[30] (
	.clk(clk_clk),
	.d(\M_dc_st_data[30]~26_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[30]~q ),
	.prn(vcc));
defparam \A_dc_st_data[30] .is_wysiwyg = "true";
defparam \A_dc_st_data[30] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[30]~30 (
	.dataa(!\M_dc_st_data[30]~26_combout ),
	.datab(!\A_dc_st_data[30]~q ),
	.datac(!\d_readdata_d1[30]~q ),
	.datad(!\A_st_data[30]~q ),
	.datae(!\dc_data_wr_port_data[25]~10_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[30]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[30]~30 .extended_lut = "off";
defparam \dc_data_wr_port_data[30]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[30]~30 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[5]~27 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\M_st_data[5]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[5]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[5]~27 .extended_lut = "off";
defparam \M_dc_st_data[5]~27 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[5]~27 .shared_arith = "off";

dffeas \A_dc_st_data[5] (
	.clk(clk_clk),
	.d(\M_dc_st_data[5]~27_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[5]~q ),
	.prn(vcc));
defparam \A_dc_st_data[5] .is_wysiwyg = "true";
defparam \A_dc_st_data[5] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[5]~31 (
	.dataa(!\M_dc_st_data[5]~27_combout ),
	.datab(!\A_dc_st_data[5]~q ),
	.datac(!\d_readdata_d1[5]~q ),
	.datad(!\A_st_data[5]~q ),
	.datae(!\dc_data_wr_port_data[1]~23_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[5]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[5]~31 .extended_lut = "off";
defparam \dc_data_wr_port_data[5]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[5]~31 .shared_arith = "off";

dffeas \i_readdata_d1[10] (
	.clk(clk_clk),
	.d(i_readdata[10]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[10]~q ),
	.prn(vcc));
defparam \i_readdata_d1[10] .is_wysiwyg = "true";
defparam \i_readdata_d1[10] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[4]~28 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\M_st_data[4]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[4]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[4]~28 .extended_lut = "off";
defparam \M_dc_st_data[4]~28 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[4]~28 .shared_arith = "off";

dffeas \A_dc_st_data[4] (
	.clk(clk_clk),
	.d(\M_dc_st_data[4]~28_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[4]~q ),
	.prn(vcc));
defparam \A_dc_st_data[4] .is_wysiwyg = "true";
defparam \A_dc_st_data[4] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[4]~32 (
	.dataa(!\M_dc_st_data[4]~28_combout ),
	.datab(!\A_dc_st_data[4]~q ),
	.datac(!\d_readdata_d1[4]~q ),
	.datad(!\A_st_data[4]~q ),
	.datae(!\dc_data_wr_port_data[1]~23_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[4]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[4]~32 .extended_lut = "off";
defparam \dc_data_wr_port_data[4]~32 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[4]~32 .shared_arith = "off";

dffeas \i_readdata_d1[9] (
	.clk(clk_clk),
	.d(i_readdata[9]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[9]~q ),
	.prn(vcc));
defparam \i_readdata_d1[9] .is_wysiwyg = "true";
defparam \i_readdata_d1[9] .power_up = "low";

cyclonev_lcell_comb \M_dc_st_data[3]~29 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\M_st_data[3]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[3]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[3]~29 .extended_lut = "off";
defparam \M_dc_st_data[3]~29 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[3]~29 .shared_arith = "off";

dffeas \A_dc_st_data[3] (
	.clk(clk_clk),
	.d(\M_dc_st_data[3]~29_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[3]~q ),
	.prn(vcc));
defparam \A_dc_st_data[3] .is_wysiwyg = "true";
defparam \A_dc_st_data[3] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[3]~33 (
	.dataa(!\M_dc_st_data[3]~29_combout ),
	.datab(!\A_dc_st_data[3]~q ),
	.datac(!\d_readdata_d1[3]~q ),
	.datad(!\A_st_data[3]~q ),
	.datae(!\dc_data_wr_port_data[1]~23_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[3]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[3]~33 .extended_lut = "off";
defparam \dc_data_wr_port_data[3]~33 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[3]~33 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[1]~30 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\M_st_data[1]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[1]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[1]~30 .extended_lut = "off";
defparam \M_dc_st_data[1]~30 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[1]~30 .shared_arith = "off";

dffeas \A_dc_st_data[1] (
	.clk(clk_clk),
	.d(\M_dc_st_data[1]~30_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[1]~q ),
	.prn(vcc));
defparam \A_dc_st_data[1] .is_wysiwyg = "true";
defparam \A_dc_st_data[1] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[1]~34 (
	.dataa(!\M_dc_st_data[1]~30_combout ),
	.datab(!\A_dc_st_data[1]~q ),
	.datac(!\d_readdata_d1[1]~q ),
	.datad(!\A_st_data[1]~q ),
	.datae(!\dc_data_wr_port_data[1]~23_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[1]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[1]~34 .extended_lut = "off";
defparam \dc_data_wr_port_data[1]~34 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[1]~34 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_st_data[0]~31 (
	.dataa(!\M_mem_byte_en[0]~q ),
	.datab(!\M_st_data[0]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_st_data[0]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_st_data[0]~31 .extended_lut = "off";
defparam \M_dc_st_data[0]~31 .lut_mask = 64'h2727272727272727;
defparam \M_dc_st_data[0]~31 .shared_arith = "off";

dffeas \A_dc_st_data[0] (
	.clk(clk_clk),
	.d(\M_dc_st_data[0]~31_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_st_data[0]~q ),
	.prn(vcc));
defparam \A_dc_st_data[0] .is_wysiwyg = "true";
defparam \A_dc_st_data[0] .power_up = "low";

cyclonev_lcell_comb \dc_data_wr_port_data[0]~35 (
	.dataa(!\M_dc_st_data[0]~31_combout ),
	.datab(!\A_dc_st_data[0]~q ),
	.datac(!\d_readdata_d1[0]~q ),
	.datad(!\A_st_data[0]~q ),
	.datae(!\dc_data_wr_port_data[1]~23_combout ),
	.dataf(!\A_dc_fill_active~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\dc_data_wr_port_data[0]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \dc_data_wr_port_data[0]~35 .extended_lut = "off";
defparam \dc_data_wr_port_data[0]~35 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \dc_data_wr_port_data[0]~35 .shared_arith = "off";

dffeas \A_dc_rd_data[6] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[6]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[6] .is_wysiwyg = "true";
defparam \A_dc_rd_data[6] .power_up = "low";

dffeas \A_dc_rd_data[4] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[4]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[4] .is_wysiwyg = "true";
defparam \A_dc_rd_data[4] .power_up = "low";

dffeas \A_dc_rd_data[7] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[7]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[7] .is_wysiwyg = "true";
defparam \A_dc_rd_data[7] .power_up = "low";

dffeas \A_dc_rd_data[5] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[5]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[5] .is_wysiwyg = "true";
defparam \A_dc_rd_data[5] .power_up = "low";

dffeas \i_readdata_d1[21] (
	.clk(clk_clk),
	.d(i_readdata[21]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[21]~q ),
	.prn(vcc));
defparam \i_readdata_d1[21] .is_wysiwyg = "true";
defparam \i_readdata_d1[21] .power_up = "low";

dffeas \i_readdata_d1[20] (
	.clk(clk_clk),
	.d(i_readdata[20]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[20]~q ),
	.prn(vcc));
defparam \i_readdata_d1[20] .is_wysiwyg = "true";
defparam \i_readdata_d1[20] .power_up = "low";

dffeas clr_break_line(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\clr_break_line~q ),
	.prn(vcc));
defparam clr_break_line.is_wysiwyg = "true";
defparam clr_break_line.power_up = "low";

cyclonev_lcell_comb ic_tag_clr_valid_bits_nxt(
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\clr_break_line~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_clr_valid_bits_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_tag_clr_valid_bits_nxt.extended_lut = "off";
defparam ic_tag_clr_valid_bits_nxt.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam ic_tag_clr_valid_bits_nxt.shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~7 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_crst~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~7 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~7 .lut_mask = 64'h7777777777777777;
defparam \ic_tag_wraddress_nxt~7 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[0]~8 (
	.dataa(!\M_alu_result[5]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~3_combout ),
	.datad(!\clr_break_line~q ),
	.datae(!\ic_tag_wraddress_nxt~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[0]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[0]~8 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[0]~8 .lut_mask = 64'hFF7FDF5FFF7FDF5F;
defparam \ic_tag_wraddress_nxt[0]~8 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[1]~9 (
	.dataa(!\clr_break_line~q ),
	.datab(!\ic_tag_wraddress_nxt~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[1]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[1]~9 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[1]~9 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \ic_tag_wraddress_nxt[1]~9 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[1]~10 (
	.dataa(!\M_alu_result[6]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~2_combout ),
	.datad(!\ic_tag_wraddress_nxt[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[1]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[1]~10 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[1]~10 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \ic_tag_wraddress_nxt[1]~10 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[2]~11 (
	.dataa(!\M_alu_result[7]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~6_combout ),
	.datad(!\ic_tag_wraddress_nxt[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[2]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[2]~11 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[2]~11 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \ic_tag_wraddress_nxt[2]~11 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[3]~12 (
	.dataa(!\M_alu_result[8]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~5_combout ),
	.datad(!\ic_tag_wraddress_nxt[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[3]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[3]~12 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[3]~12 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \ic_tag_wraddress_nxt[3]~12 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[4]~13 (
	.dataa(!\M_alu_result[9]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~4_combout ),
	.datad(!\ic_tag_wraddress_nxt[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[4]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[4]~13 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[4]~13 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \ic_tag_wraddress_nxt[4]~13 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[5]~14 (
	.dataa(!\M_alu_result[10]~q ),
	.datab(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datac(!\ic_tag_wraddress_nxt~1_combout ),
	.datad(!\ic_tag_wraddress_nxt[1]~9_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[5]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[5]~14 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[5]~14 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \ic_tag_wraddress_nxt[5]~14 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt[6]~15 (
	.dataa(!\M_alu_result[11]~q ),
	.datab(!\ic_tag_wraddress_nxt~0_combout ),
	.datac(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datad(!\clr_break_line~q ),
	.datae(!\ic_tag_wraddress_nxt~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt[6]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt[6]~15 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt[6]~15 .lut_mask = 64'hFF7FF777FF7FF777;
defparam \ic_tag_wraddress_nxt[6]~15 .shared_arith = "off";

dffeas \i_readdata_d1[7] (
	.clk(clk_clk),
	.d(i_readdata[7]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[7]~q ),
	.prn(vcc));
defparam \i_readdata_d1[7] .is_wysiwyg = "true";
defparam \i_readdata_d1[7] .power_up = "low";

dffeas \i_readdata_d1[6] (
	.clk(clk_clk),
	.d(i_readdata[6]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdata_d1[6]~q ),
	.prn(vcc));
defparam \i_readdata_d1[6] .is_wysiwyg = "true";
defparam \i_readdata_d1[6] .power_up = "low";

dffeas \E_bht_data[0] (
	.clk(clk_clk),
	.d(\D_bht_data[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_data[0]~q ),
	.prn(vcc));
defparam \E_bht_data[0] .is_wysiwyg = "true";
defparam \E_bht_data[0] .power_up = "low";

cyclonev_lcell_comb E_br_mispredict(
	.dataa(!\E_valid~1_combout ),
	.datab(!\E_bht_data[1]~q ),
	.datac(!\Add17~61_sumout ),
	.datad(!\E_br_result~0_combout ),
	.datae(!\E_br_result~1_combout ),
	.dataf(!\E_ctrl_br_cond~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_mispredict~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_br_mispredict.extended_lut = "off";
defparam E_br_mispredict.lut_mask = 64'h7DD7D77DFFFFFFFF;
defparam E_br_mispredict.shared_arith = "off";

dffeas \E_bht_ptr[0] (
	.clk(clk_clk),
	.d(\D_bht_ptr[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[0]~q ),
	.prn(vcc));
defparam \E_bht_ptr[0] .is_wysiwyg = "true";
defparam \E_bht_ptr[0] .power_up = "low";

dffeas \E_bht_ptr[1] (
	.clk(clk_clk),
	.d(\D_bht_ptr[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[1]~q ),
	.prn(vcc));
defparam \E_bht_ptr[1] .is_wysiwyg = "true";
defparam \E_bht_ptr[1] .power_up = "low";

dffeas \E_bht_ptr[2] (
	.clk(clk_clk),
	.d(\D_bht_ptr[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[2]~q ),
	.prn(vcc));
defparam \E_bht_ptr[2] .is_wysiwyg = "true";
defparam \E_bht_ptr[2] .power_up = "low";

dffeas \E_bht_ptr[3] (
	.clk(clk_clk),
	.d(\D_bht_ptr[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[3]~q ),
	.prn(vcc));
defparam \E_bht_ptr[3] .is_wysiwyg = "true";
defparam \E_bht_ptr[3] .power_up = "low";

dffeas \E_bht_ptr[4] (
	.clk(clk_clk),
	.d(\D_bht_ptr[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[4]~q ),
	.prn(vcc));
defparam \E_bht_ptr[4] .is_wysiwyg = "true";
defparam \E_bht_ptr[4] .power_up = "low";

dffeas \E_bht_ptr[5] (
	.clk(clk_clk),
	.d(\D_bht_ptr[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[5]~q ),
	.prn(vcc));
defparam \E_bht_ptr[5] .is_wysiwyg = "true";
defparam \E_bht_ptr[5] .power_up = "low";

dffeas \E_bht_ptr[6] (
	.clk(clk_clk),
	.d(\D_bht_ptr[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[6]~q ),
	.prn(vcc));
defparam \E_bht_ptr[6] .is_wysiwyg = "true";
defparam \E_bht_ptr[6] .power_up = "low";

dffeas \E_bht_ptr[7] (
	.clk(clk_clk),
	.d(\D_bht_ptr[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_ptr[7]~q ),
	.prn(vcc));
defparam \E_bht_ptr[7] .is_wysiwyg = "true";
defparam \E_bht_ptr[7] .power_up = "low";

cyclonev_lcell_comb \M_br_cond_taken_history[0]~0 (
	.dataa(!\A_mem_stall~q ),
	.datab(!\A_mul_stall~q ),
	.datac(!\E_ctrl_br_cond~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_br_cond_taken_history[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_br_cond_taken_history[0]~0 .extended_lut = "off";
defparam \M_br_cond_taken_history[0]~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \M_br_cond_taken_history[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \M_br_cond_taken_history[0]~1 (
	.dataa(!\E_valid~0_combout ),
	.datab(!\E_hbreak_req~0_combout ),
	.datac(!\Equal209~0_combout ),
	.datad(!\E_hbreak_req~1_combout ),
	.datae(!\hbreak_req~0_combout ),
	.dataf(!\M_br_cond_taken_history[0]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_br_cond_taken_history[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_br_cond_taken_history[0]~1 .extended_lut = "off";
defparam \M_br_cond_taken_history[0]~1 .lut_mask = 64'hFFFF7FFFFFFFFFFF;
defparam \M_br_cond_taken_history[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~0 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~0 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \ic_fill_valid_bits_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb ic_fill_valid_bits_en(
	.dataa(!\ic_fill_dp_offset_en~0_combout ),
	.datab(!\ic_tag_clr_valid_bits_nxt~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_en~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_fill_valid_bits_en.extended_lut = "off";
defparam ic_fill_valid_bits_en.lut_mask = 64'h7777777777777777;
defparam ic_fill_valid_bits_en.shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~1 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~1 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~1 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \ic_fill_valid_bits_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~2 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~2 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~2 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \ic_fill_valid_bits_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~3 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~3 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~3 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \ic_fill_valid_bits_nxt~3 .shared_arith = "off";

dffeas \D_bht_data[0] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_data[0]~q ),
	.prn(vcc));
defparam \D_bht_data[0] .is_wysiwyg = "true";
defparam \D_bht_data[0] .power_up = "low";

dffeas \D_bht_ptr[0] (
	.clk(clk_clk),
	.d(\F_bht_ptr[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[0]~q ),
	.prn(vcc));
defparam \D_bht_ptr[0] .is_wysiwyg = "true";
defparam \D_bht_ptr[0] .power_up = "low";

dffeas \D_bht_ptr[1] (
	.clk(clk_clk),
	.d(\F_bht_ptr[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[1]~q ),
	.prn(vcc));
defparam \D_bht_ptr[1] .is_wysiwyg = "true";
defparam \D_bht_ptr[1] .power_up = "low";

dffeas \D_bht_ptr[2] (
	.clk(clk_clk),
	.d(\F_bht_ptr[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[2]~q ),
	.prn(vcc));
defparam \D_bht_ptr[2] .is_wysiwyg = "true";
defparam \D_bht_ptr[2] .power_up = "low";

dffeas \D_bht_ptr[3] (
	.clk(clk_clk),
	.d(\F_bht_ptr[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[3]~q ),
	.prn(vcc));
defparam \D_bht_ptr[3] .is_wysiwyg = "true";
defparam \D_bht_ptr[3] .power_up = "low";

dffeas \D_bht_ptr[4] (
	.clk(clk_clk),
	.d(\F_bht_ptr[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[4]~q ),
	.prn(vcc));
defparam \D_bht_ptr[4] .is_wysiwyg = "true";
defparam \D_bht_ptr[4] .power_up = "low";

dffeas \D_bht_ptr[5] (
	.clk(clk_clk),
	.d(\F_bht_ptr[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[5]~q ),
	.prn(vcc));
defparam \D_bht_ptr[5] .is_wysiwyg = "true";
defparam \D_bht_ptr[5] .power_up = "low";

dffeas \D_bht_ptr[6] (
	.clk(clk_clk),
	.d(\F_bht_ptr[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[6]~q ),
	.prn(vcc));
defparam \D_bht_ptr[6] .is_wysiwyg = "true";
defparam \D_bht_ptr[6] .power_up = "low";

dffeas \D_bht_ptr[7] (
	.clk(clk_clk),
	.d(\F_bht_ptr[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_ptr[7]~q ),
	.prn(vcc));
defparam \D_bht_ptr[7] .is_wysiwyg = "true";
defparam \D_bht_ptr[7] .power_up = "low";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~4 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~4 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~4 .lut_mask = 64'hFFFBFFFFFFFBFFFF;
defparam \ic_fill_valid_bits_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~5 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~5 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~5 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \ic_fill_valid_bits_nxt~5 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~6 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~6 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~6 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \ic_fill_valid_bits_nxt~6 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_valid_bits_nxt~7 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datac(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_valid_bits[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_valid_bits_nxt~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_valid_bits_nxt~7 .extended_lut = "off";
defparam \ic_fill_valid_bits_nxt~7 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \ic_fill_valid_bits_nxt~7 .shared_arith = "off";

dffeas \M_src2[0] (
	.clk(clk_clk),
	.d(\E_src2[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[0]~q ),
	.prn(vcc));
defparam \M_src2[0] .is_wysiwyg = "true";
defparam \M_src2[0] .power_up = "low";

dffeas \M_src2[1] (
	.clk(clk_clk),
	.d(\E_src2[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[1]~q ),
	.prn(vcc));
defparam \M_src2[1] .is_wysiwyg = "true";
defparam \M_src2[1] .power_up = "low";

dffeas \M_src2[2] (
	.clk(clk_clk),
	.d(\E_src2[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[2]~q ),
	.prn(vcc));
defparam \M_src2[2] .is_wysiwyg = "true";
defparam \M_src2[2] .power_up = "low";

dffeas \M_src2[3] (
	.clk(clk_clk),
	.d(\E_src2[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[3]~q ),
	.prn(vcc));
defparam \M_src2[3] .is_wysiwyg = "true";
defparam \M_src2[3] .power_up = "low";

dffeas \M_src2[4] (
	.clk(clk_clk),
	.d(\E_src2[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[4]~q ),
	.prn(vcc));
defparam \M_src2[4] .is_wysiwyg = "true";
defparam \M_src2[4] .power_up = "low";

dffeas \M_src2[5] (
	.clk(clk_clk),
	.d(\E_src2[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[5]~q ),
	.prn(vcc));
defparam \M_src2[5] .is_wysiwyg = "true";
defparam \M_src2[5] .power_up = "low";

dffeas \M_src2[6] (
	.clk(clk_clk),
	.d(\E_src2[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[6]~q ),
	.prn(vcc));
defparam \M_src2[6] .is_wysiwyg = "true";
defparam \M_src2[6] .power_up = "low";

dffeas \M_src2[7] (
	.clk(clk_clk),
	.d(\E_src2[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[7]~q ),
	.prn(vcc));
defparam \M_src2[7] .is_wysiwyg = "true";
defparam \M_src2[7] .power_up = "low";

dffeas \M_src2[8] (
	.clk(clk_clk),
	.d(\E_src2[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[8]~q ),
	.prn(vcc));
defparam \M_src2[8] .is_wysiwyg = "true";
defparam \M_src2[8] .power_up = "low";

dffeas \M_src2[9] (
	.clk(clk_clk),
	.d(\E_src2[9]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[9]~q ),
	.prn(vcc));
defparam \M_src2[9] .is_wysiwyg = "true";
defparam \M_src2[9] .power_up = "low";

dffeas \M_src2[10] (
	.clk(clk_clk),
	.d(\E_src2[10]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[10]~q ),
	.prn(vcc));
defparam \M_src2[10] .is_wysiwyg = "true";
defparam \M_src2[10] .power_up = "low";

dffeas \M_src2[11] (
	.clk(clk_clk),
	.d(\E_src2[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[11]~q ),
	.prn(vcc));
defparam \M_src2[11] .is_wysiwyg = "true";
defparam \M_src2[11] .power_up = "low";

dffeas \M_src2[12] (
	.clk(clk_clk),
	.d(\E_src2[12]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[12]~q ),
	.prn(vcc));
defparam \M_src2[12] .is_wysiwyg = "true";
defparam \M_src2[12] .power_up = "low";

dffeas \M_src2[13] (
	.clk(clk_clk),
	.d(\E_src2[13]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[13]~q ),
	.prn(vcc));
defparam \M_src2[13] .is_wysiwyg = "true";
defparam \M_src2[13] .power_up = "low";

dffeas \M_src2[14] (
	.clk(clk_clk),
	.d(\E_src2[14]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[14]~q ),
	.prn(vcc));
defparam \M_src2[14] .is_wysiwyg = "true";
defparam \M_src2[14] .power_up = "low";

dffeas \M_src2[15] (
	.clk(clk_clk),
	.d(\E_src2[15]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[15]~q ),
	.prn(vcc));
defparam \M_src2[15] .is_wysiwyg = "true";
defparam \M_src2[15] .power_up = "low";

dffeas \M_src1[0] (
	.clk(clk_clk),
	.d(\E_src1[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[0]~q ),
	.prn(vcc));
defparam \M_src1[0] .is_wysiwyg = "true";
defparam \M_src1[0] .power_up = "low";

dffeas \M_src1[1] (
	.clk(clk_clk),
	.d(\E_src1[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[1]~q ),
	.prn(vcc));
defparam \M_src1[1] .is_wysiwyg = "true";
defparam \M_src1[1] .power_up = "low";

dffeas \M_src1[2] (
	.clk(clk_clk),
	.d(\E_src1[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[2]~q ),
	.prn(vcc));
defparam \M_src1[2] .is_wysiwyg = "true";
defparam \M_src1[2] .power_up = "low";

dffeas \M_src1[3] (
	.clk(clk_clk),
	.d(\E_src1[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[3]~q ),
	.prn(vcc));
defparam \M_src1[3] .is_wysiwyg = "true";
defparam \M_src1[3] .power_up = "low";

dffeas \M_src1[4] (
	.clk(clk_clk),
	.d(\E_src1[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[4]~q ),
	.prn(vcc));
defparam \M_src1[4] .is_wysiwyg = "true";
defparam \M_src1[4] .power_up = "low";

dffeas \M_src1[5] (
	.clk(clk_clk),
	.d(\E_src1[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[5]~q ),
	.prn(vcc));
defparam \M_src1[5] .is_wysiwyg = "true";
defparam \M_src1[5] .power_up = "low";

dffeas \M_src1[6] (
	.clk(clk_clk),
	.d(\E_src1[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[6]~q ),
	.prn(vcc));
defparam \M_src1[6] .is_wysiwyg = "true";
defparam \M_src1[6] .power_up = "low";

dffeas \M_src1[7] (
	.clk(clk_clk),
	.d(\E_src1[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[7]~q ),
	.prn(vcc));
defparam \M_src1[7] .is_wysiwyg = "true";
defparam \M_src1[7] .power_up = "low";

dffeas \M_src1[8] (
	.clk(clk_clk),
	.d(\E_src1[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[8]~q ),
	.prn(vcc));
defparam \M_src1[8] .is_wysiwyg = "true";
defparam \M_src1[8] .power_up = "low";

dffeas \M_src1[9] (
	.clk(clk_clk),
	.d(\E_src1[9]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[9]~q ),
	.prn(vcc));
defparam \M_src1[9] .is_wysiwyg = "true";
defparam \M_src1[9] .power_up = "low";

dffeas \M_src1[10] (
	.clk(clk_clk),
	.d(\E_src1[10]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[10]~q ),
	.prn(vcc));
defparam \M_src1[10] .is_wysiwyg = "true";
defparam \M_src1[10] .power_up = "low";

dffeas \M_src1[11] (
	.clk(clk_clk),
	.d(\E_src1[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[11]~q ),
	.prn(vcc));
defparam \M_src1[11] .is_wysiwyg = "true";
defparam \M_src1[11] .power_up = "low";

dffeas \M_src1[12] (
	.clk(clk_clk),
	.d(\E_src1[12]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[12]~q ),
	.prn(vcc));
defparam \M_src1[12] .is_wysiwyg = "true";
defparam \M_src1[12] .power_up = "low";

dffeas \M_src1[13] (
	.clk(clk_clk),
	.d(\E_src1[13]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[13]~q ),
	.prn(vcc));
defparam \M_src1[13] .is_wysiwyg = "true";
defparam \M_src1[13] .power_up = "low";

dffeas \M_src1[14] (
	.clk(clk_clk),
	.d(\E_src1[14]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[14]~q ),
	.prn(vcc));
defparam \M_src1[14] .is_wysiwyg = "true";
defparam \M_src1[14] .power_up = "low";

dffeas \M_src1[15] (
	.clk(clk_clk),
	.d(\E_src1[15]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[15]~q ),
	.prn(vcc));
defparam \M_src1[15] .is_wysiwyg = "true";
defparam \M_src1[15] .power_up = "low";

dffeas \F_bht_ptr[0] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[0]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[0]~q ),
	.prn(vcc));
defparam \F_bht_ptr[0] .is_wysiwyg = "true";
defparam \F_bht_ptr[0] .power_up = "low";

dffeas \F_bht_ptr[1] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[1]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[1]~q ),
	.prn(vcc));
defparam \F_bht_ptr[1] .is_wysiwyg = "true";
defparam \F_bht_ptr[1] .power_up = "low";

dffeas \F_bht_ptr[2] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[2]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[2]~q ),
	.prn(vcc));
defparam \F_bht_ptr[2] .is_wysiwyg = "true";
defparam \F_bht_ptr[2] .power_up = "low";

dffeas \F_bht_ptr[3] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[3]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[3]~q ),
	.prn(vcc));
defparam \F_bht_ptr[3] .is_wysiwyg = "true";
defparam \F_bht_ptr[3] .power_up = "low";

dffeas \F_bht_ptr[4] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[4]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[4]~q ),
	.prn(vcc));
defparam \F_bht_ptr[4] .is_wysiwyg = "true";
defparam \F_bht_ptr[4] .power_up = "low";

dffeas \F_bht_ptr[5] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[5]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[5]~q ),
	.prn(vcc));
defparam \F_bht_ptr[5] .is_wysiwyg = "true";
defparam \F_bht_ptr[5] .power_up = "low";

dffeas \F_bht_ptr[6] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[6]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[6]~q ),
	.prn(vcc));
defparam \F_bht_ptr[6] .is_wysiwyg = "true";
defparam \F_bht_ptr[6] .power_up = "low";

dffeas \F_bht_ptr[7] (
	.clk(clk_clk),
	.d(\F_bht_ptr_nxt[7]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_bht_ptr[7]~q ),
	.prn(vcc));
defparam \F_bht_ptr[7] .is_wysiwyg = "true";
defparam \F_bht_ptr[7] .power_up = "low";

dffeas \M_src2[16] (
	.clk(clk_clk),
	.d(\E_src2[16]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[16]~q ),
	.prn(vcc));
defparam \M_src2[16] .is_wysiwyg = "true";
defparam \M_src2[16] .power_up = "low";

dffeas \M_src2[17] (
	.clk(clk_clk),
	.d(\E_src2[17]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[17]~q ),
	.prn(vcc));
defparam \M_src2[17] .is_wysiwyg = "true";
defparam \M_src2[17] .power_up = "low";

dffeas \M_src2[18] (
	.clk(clk_clk),
	.d(\E_src2[18]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[18]~q ),
	.prn(vcc));
defparam \M_src2[18] .is_wysiwyg = "true";
defparam \M_src2[18] .power_up = "low";

dffeas \M_src2[19] (
	.clk(clk_clk),
	.d(\E_src2[19]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[19]~q ),
	.prn(vcc));
defparam \M_src2[19] .is_wysiwyg = "true";
defparam \M_src2[19] .power_up = "low";

dffeas \M_src2[20] (
	.clk(clk_clk),
	.d(\E_src2[20]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[20]~q ),
	.prn(vcc));
defparam \M_src2[20] .is_wysiwyg = "true";
defparam \M_src2[20] .power_up = "low";

dffeas \M_src2[21] (
	.clk(clk_clk),
	.d(\E_src2[21]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[21]~q ),
	.prn(vcc));
defparam \M_src2[21] .is_wysiwyg = "true";
defparam \M_src2[21] .power_up = "low";

dffeas \M_src2[22] (
	.clk(clk_clk),
	.d(\E_src2[22]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[22]~q ),
	.prn(vcc));
defparam \M_src2[22] .is_wysiwyg = "true";
defparam \M_src2[22] .power_up = "low";

dffeas \M_src2[23] (
	.clk(clk_clk),
	.d(\E_src2[23]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[23]~q ),
	.prn(vcc));
defparam \M_src2[23] .is_wysiwyg = "true";
defparam \M_src2[23] .power_up = "low";

dffeas \M_src2[24] (
	.clk(clk_clk),
	.d(\E_src2[24]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[24]~q ),
	.prn(vcc));
defparam \M_src2[24] .is_wysiwyg = "true";
defparam \M_src2[24] .power_up = "low";

dffeas \M_src2[25] (
	.clk(clk_clk),
	.d(\E_src2[25]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[25]~q ),
	.prn(vcc));
defparam \M_src2[25] .is_wysiwyg = "true";
defparam \M_src2[25] .power_up = "low";

dffeas \M_src2[26] (
	.clk(clk_clk),
	.d(\E_src2[26]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[26]~q ),
	.prn(vcc));
defparam \M_src2[26] .is_wysiwyg = "true";
defparam \M_src2[26] .power_up = "low";

dffeas \M_src2[27] (
	.clk(clk_clk),
	.d(\E_src2[27]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[27]~q ),
	.prn(vcc));
defparam \M_src2[27] .is_wysiwyg = "true";
defparam \M_src2[27] .power_up = "low";

dffeas \M_src2[28] (
	.clk(clk_clk),
	.d(\E_src2[28]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[28]~q ),
	.prn(vcc));
defparam \M_src2[28] .is_wysiwyg = "true";
defparam \M_src2[28] .power_up = "low";

dffeas \M_src2[29] (
	.clk(clk_clk),
	.d(\E_src2[29]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[29]~q ),
	.prn(vcc));
defparam \M_src2[29] .is_wysiwyg = "true";
defparam \M_src2[29] .power_up = "low";

dffeas \M_src2[30] (
	.clk(clk_clk),
	.d(\E_src2[30]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[30]~q ),
	.prn(vcc));
defparam \M_src2[30] .is_wysiwyg = "true";
defparam \M_src2[30] .power_up = "low";

dffeas \M_src2[31] (
	.clk(clk_clk),
	.d(\E_src2[31]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src2[31]~q ),
	.prn(vcc));
defparam \M_src2[31] .is_wysiwyg = "true";
defparam \M_src2[31] .power_up = "low";

dffeas \A_dc_rd_data[31] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[31]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[31] .is_wysiwyg = "true";
defparam \A_dc_rd_data[31] .power_up = "low";

dffeas \A_dc_rd_data[29] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[29]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[29] .is_wysiwyg = "true";
defparam \A_dc_rd_data[29] .power_up = "low";

dffeas \A_dc_rd_data[28] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[28]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[28] .is_wysiwyg = "true";
defparam \A_dc_rd_data[28] .power_up = "low";

dffeas \A_dc_rd_data[30] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_rd_data[30]~q ),
	.prn(vcc));
defparam \A_dc_rd_data[30] .is_wysiwyg = "true";
defparam \A_dc_rd_data[30] .power_up = "low";

dffeas \M_src1[16] (
	.clk(clk_clk),
	.d(\E_src1[16]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[16]~q ),
	.prn(vcc));
defparam \M_src1[16] .is_wysiwyg = "true";
defparam \M_src1[16] .power_up = "low";

dffeas \M_src1[17] (
	.clk(clk_clk),
	.d(\E_src1[17]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[17]~q ),
	.prn(vcc));
defparam \M_src1[17] .is_wysiwyg = "true";
defparam \M_src1[17] .power_up = "low";

dffeas \M_src1[18] (
	.clk(clk_clk),
	.d(\E_src1[18]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[18]~q ),
	.prn(vcc));
defparam \M_src1[18] .is_wysiwyg = "true";
defparam \M_src1[18] .power_up = "low";

dffeas \M_src1[19] (
	.clk(clk_clk),
	.d(\E_src1[19]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[19]~q ),
	.prn(vcc));
defparam \M_src1[19] .is_wysiwyg = "true";
defparam \M_src1[19] .power_up = "low";

dffeas \M_src1[20] (
	.clk(clk_clk),
	.d(\E_src1[20]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[20]~q ),
	.prn(vcc));
defparam \M_src1[20] .is_wysiwyg = "true";
defparam \M_src1[20] .power_up = "low";

dffeas \M_src1[21] (
	.clk(clk_clk),
	.d(\E_src1[21]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[21]~q ),
	.prn(vcc));
defparam \M_src1[21] .is_wysiwyg = "true";
defparam \M_src1[21] .power_up = "low";

dffeas \M_src1[22] (
	.clk(clk_clk),
	.d(\E_src1[22]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[22]~q ),
	.prn(vcc));
defparam \M_src1[22] .is_wysiwyg = "true";
defparam \M_src1[22] .power_up = "low";

dffeas \M_src1[23] (
	.clk(clk_clk),
	.d(\E_src1[23]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[23]~q ),
	.prn(vcc));
defparam \M_src1[23] .is_wysiwyg = "true";
defparam \M_src1[23] .power_up = "low";

dffeas \M_src1[24] (
	.clk(clk_clk),
	.d(\E_src1[24]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[24]~q ),
	.prn(vcc));
defparam \M_src1[24] .is_wysiwyg = "true";
defparam \M_src1[24] .power_up = "low";

dffeas \M_src1[25] (
	.clk(clk_clk),
	.d(\E_src1[25]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[25]~q ),
	.prn(vcc));
defparam \M_src1[25] .is_wysiwyg = "true";
defparam \M_src1[25] .power_up = "low";

dffeas \M_src1[26] (
	.clk(clk_clk),
	.d(\E_src1[26]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[26]~q ),
	.prn(vcc));
defparam \M_src1[26] .is_wysiwyg = "true";
defparam \M_src1[26] .power_up = "low";

dffeas \M_src1[27] (
	.clk(clk_clk),
	.d(\E_src1[27]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[27]~q ),
	.prn(vcc));
defparam \M_src1[27] .is_wysiwyg = "true";
defparam \M_src1[27] .power_up = "low";

dffeas \M_src1[28] (
	.clk(clk_clk),
	.d(\E_src1[28]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[28]~q ),
	.prn(vcc));
defparam \M_src1[28] .is_wysiwyg = "true";
defparam \M_src1[28] .power_up = "low";

dffeas \M_src1[29] (
	.clk(clk_clk),
	.d(\E_src1[29]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[29]~q ),
	.prn(vcc));
defparam \M_src1[29] .is_wysiwyg = "true";
defparam \M_src1[29] .power_up = "low";

dffeas \M_src1[30] (
	.clk(clk_clk),
	.d(\E_src1[30]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[30]~q ),
	.prn(vcc));
defparam \M_src1[30] .is_wysiwyg = "true";
defparam \M_src1[30] .power_up = "low";

dffeas \M_src1[31] (
	.clk(clk_clk),
	.d(\E_src1[31]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_src1[31]~q ),
	.prn(vcc));
defparam \M_src1[31] .is_wysiwyg = "true";
defparam \M_src1[31] .power_up = "low";

cyclonev_lcell_comb \ic_tag_clr_valid_bits~0 (
	.dataa(!\ic_tag_clr_valid_bits_nxt~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_clr_valid_bits~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_clr_valid_bits~0 .extended_lut = "off";
defparam \ic_tag_clr_valid_bits~0 .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \ic_tag_clr_valid_bits~0 .shared_arith = "off";

cyclonev_lcell_comb \M_br_mispredict~_wirecell (
	.dataa(!\M_br_mispredict~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_br_mispredict~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_br_mispredict~_wirecell .extended_lut = "off";
defparam \M_br_mispredict~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \M_br_mispredict~_wirecell .shared_arith = "off";

dffeas \d_address_offset_field[0] (
	.clk(clk_clk),
	.d(\d_address_offset_field_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_address_offset_field[1]~3_combout ),
	.q(d_address_offset_field_0),
	.prn(vcc));
defparam \d_address_offset_field[0] .is_wysiwyg = "true";
defparam \d_address_offset_field[0] .power_up = "low";

dffeas \d_write~reg0 (
	.clk(clk_clk),
	.d(\d_write_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_write),
	.prn(vcc));
defparam \d_write~reg0 .is_wysiwyg = "true";
defparam \d_write~reg0 .power_up = "low";

dffeas \d_address_tag_field[2] (
	.clk(clk_clk),
	.d(\d_address_tag_field_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_tag_field_2),
	.prn(vcc));
defparam \d_address_tag_field[2] .is_wysiwyg = "true";
defparam \d_address_tag_field[2] .power_up = "low";

dffeas \d_address_tag_field[1] (
	.clk(clk_clk),
	.d(\d_address_tag_field_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_tag_field_1),
	.prn(vcc));
defparam \d_address_tag_field[1] .is_wysiwyg = "true";
defparam \d_address_tag_field[1] .power_up = "low";

dffeas \d_address_tag_field[0] (
	.clk(clk_clk),
	.d(\d_address_tag_field_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_tag_field_0),
	.prn(vcc));
defparam \d_address_tag_field[0] .is_wysiwyg = "true";
defparam \d_address_tag_field[0] .power_up = "low";

dffeas \d_address_line_field[5] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[5]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_5),
	.prn(vcc));
defparam \d_address_line_field[5] .is_wysiwyg = "true";
defparam \d_address_line_field[5] .power_up = "low";

dffeas \d_address_line_field[4] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[4]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_4),
	.prn(vcc));
defparam \d_address_line_field[4] .is_wysiwyg = "true";
defparam \d_address_line_field[4] .power_up = "low";

dffeas \d_address_line_field[3] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[3]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_3),
	.prn(vcc));
defparam \d_address_line_field[3] .is_wysiwyg = "true";
defparam \d_address_line_field[3] .power_up = "low";

dffeas \d_address_line_field[2] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[2]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_2),
	.prn(vcc));
defparam \d_address_line_field[2] .is_wysiwyg = "true";
defparam \d_address_line_field[2] .power_up = "low";

dffeas \d_address_line_field[1] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[1]~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_1),
	.prn(vcc));
defparam \d_address_line_field[1] .is_wysiwyg = "true";
defparam \d_address_line_field[1] .power_up = "low";

dffeas \d_address_line_field[0] (
	.clk(clk_clk),
	.d(\d_address_line_field_nxt[0]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_address_line_field_0),
	.prn(vcc));
defparam \d_address_line_field[0] .is_wysiwyg = "true";
defparam \d_address_line_field[0] .power_up = "low";

dffeas \d_address_offset_field[2] (
	.clk(clk_clk),
	.d(\d_address_offset_field_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_address_offset_field[1]~3_combout ),
	.q(d_address_offset_field_2),
	.prn(vcc));
defparam \d_address_offset_field[2] .is_wysiwyg = "true";
defparam \d_address_offset_field[2] .power_up = "low";

dffeas \d_address_offset_field[1] (
	.clk(clk_clk),
	.d(\d_address_offset_field_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_address_offset_field[1]~3_combout ),
	.q(d_address_offset_field_1),
	.prn(vcc));
defparam \d_address_offset_field[1] .is_wysiwyg = "true";
defparam \d_address_offset_field[1] .power_up = "low";

dffeas \d_writedata[11]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[11]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_11),
	.prn(vcc));
defparam \d_writedata[11]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[11]~reg0 .power_up = "low";

dffeas \d_byteenable[0]~reg0 (
	.clk(clk_clk),
	.d(\d_byteenable_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_0),
	.prn(vcc));
defparam \d_byteenable[0]~reg0 .is_wysiwyg = "true";
defparam \d_byteenable[0]~reg0 .power_up = "low";

dffeas \d_writedata[10]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[10]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_10),
	.prn(vcc));
defparam \d_writedata[10]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[10]~reg0 .power_up = "low";

dffeas \d_writedata[9]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[9]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_9),
	.prn(vcc));
defparam \d_writedata[9]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[9]~reg0 .power_up = "low";

dffeas \d_writedata[8]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[8]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_8),
	.prn(vcc));
defparam \d_writedata[8]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[8]~reg0 .power_up = "low";

dffeas \d_writedata[13]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[13]~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_13),
	.prn(vcc));
defparam \d_writedata[13]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[13]~reg0 .power_up = "low";

dffeas \d_writedata[12]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[12]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_12),
	.prn(vcc));
defparam \d_writedata[12]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[12]~reg0 .power_up = "low";

dffeas \d_writedata[21]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[21]~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_21),
	.prn(vcc));
defparam \d_writedata[21]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[21]~reg0 .power_up = "low";

dffeas \d_writedata[20]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[20]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_20),
	.prn(vcc));
defparam \d_writedata[20]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[20]~reg0 .power_up = "low";

dffeas \d_writedata[25]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[25]~8_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_25),
	.prn(vcc));
defparam \d_writedata[25]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[25]~reg0 .power_up = "low";

dffeas \d_writedata[17]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[17]~9_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_17),
	.prn(vcc));
defparam \d_writedata[17]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[17]~reg0 .power_up = "low";

dffeas \d_writedata[24]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[24]~10_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_24),
	.prn(vcc));
defparam \d_writedata[24]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[24]~reg0 .power_up = "low";

dffeas \d_writedata[16]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[16]~11_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_16),
	.prn(vcc));
defparam \d_writedata[16]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[16]~reg0 .power_up = "low";

dffeas \d_writedata[27]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[27]~12_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_27),
	.prn(vcc));
defparam \d_writedata[27]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[27]~reg0 .power_up = "low";

dffeas \d_writedata[19]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[19]~13_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_19),
	.prn(vcc));
defparam \d_writedata[19]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[19]~reg0 .power_up = "low";

dffeas \d_writedata[26]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[26]~14_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_26),
	.prn(vcc));
defparam \d_writedata[26]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[26]~reg0 .power_up = "low";

dffeas \d_writedata[18]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[18]~15_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_18),
	.prn(vcc));
defparam \d_writedata[18]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[18]~reg0 .power_up = "low";

dffeas \d_writedata[23]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[23]~16_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_23),
	.prn(vcc));
defparam \d_writedata[23]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[23]~reg0 .power_up = "low";

dffeas \d_writedata[15]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[15]~17_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_15),
	.prn(vcc));
defparam \d_writedata[15]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[15]~reg0 .power_up = "low";

dffeas \d_writedata[22]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[22]~18_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_22),
	.prn(vcc));
defparam \d_writedata[22]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[22]~reg0 .power_up = "low";

dffeas \d_writedata[14]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[14]~19_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_14),
	.prn(vcc));
defparam \d_writedata[14]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[14]~reg0 .power_up = "low";

dffeas \d_read~reg0 (
	.clk(clk_clk),
	.d(\d_read_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_read),
	.prn(vcc));
defparam \d_read~reg0 .is_wysiwyg = "true";
defparam \d_read~reg0 .power_up = "low";

dffeas \d_byteenable[1]~reg0 (
	.clk(clk_clk),
	.d(\d_byteenable_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_1),
	.prn(vcc));
defparam \d_byteenable[1]~reg0 .is_wysiwyg = "true";
defparam \d_byteenable[1]~reg0 .power_up = "low";

dffeas \d_writedata[2]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[2]~20_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_2),
	.prn(vcc));
defparam \d_writedata[2]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[2]~reg0 .power_up = "low";

dffeas \d_writedata[0]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[0]~21_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_0),
	.prn(vcc));
defparam \d_writedata[0]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[0]~reg0 .power_up = "low";

dffeas \d_writedata[3]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[3]~22_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_3),
	.prn(vcc));
defparam \d_writedata[3]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[3]~reg0 .power_up = "low";

dffeas \d_writedata[1]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[1]~23_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_1),
	.prn(vcc));
defparam \d_writedata[1]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[1]~reg0 .power_up = "low";

dffeas hbreak_enabled(
	.clk(clk_clk),
	.d(\hbreak_enabled~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always120~0_combout ),
	.q(hbreak_enabled1),
	.prn(vcc));
defparam hbreak_enabled.is_wysiwyg = "true";
defparam hbreak_enabled.power_up = "low";

dffeas \i_read~reg0 (
	.clk(clk_clk),
	.d(\i_read_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(i_read),
	.prn(vcc));
defparam \i_read~reg0 .is_wysiwyg = "true";
defparam \i_read~reg0 .power_up = "low";

dffeas \ic_fill_tag[1] (
	.clk(clk_clk),
	.d(\D_pc[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_1),
	.prn(vcc));
defparam \ic_fill_tag[1] .is_wysiwyg = "true";
defparam \ic_fill_tag[1] .power_up = "low";

dffeas \ic_fill_tag[0] (
	.clk(clk_clk),
	.d(\D_pc[10]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(ic_fill_tag_0),
	.prn(vcc));
defparam \ic_fill_tag[0] .is_wysiwyg = "true";
defparam \ic_fill_tag[0] .power_up = "low";

dffeas \ic_fill_line[6] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_6),
	.prn(vcc));
defparam \ic_fill_line[6] .is_wysiwyg = "true";
defparam \ic_fill_line[6] .power_up = "low";

dffeas \d_writedata[6]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[6]~24_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_6),
	.prn(vcc));
defparam \d_writedata[6]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[6]~reg0 .power_up = "low";

dffeas \d_writedata[4]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[4]~25_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_4),
	.prn(vcc));
defparam \d_writedata[4]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[4]~reg0 .power_up = "low";

dffeas \d_writedata[7]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[7]~26_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_7),
	.prn(vcc));
defparam \d_writedata[7]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[7]~reg0 .power_up = "low";

dffeas \d_writedata[5]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[5]~27_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_5),
	.prn(vcc));
defparam \d_writedata[5]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[5]~reg0 .power_up = "low";

dffeas \ic_fill_line[5] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_5),
	.prn(vcc));
defparam \ic_fill_line[5] .is_wysiwyg = "true";
defparam \ic_fill_line[5] .power_up = "low";

dffeas \ic_fill_ap_offset[0] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[0]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[1]~0_combout ),
	.q(ic_fill_ap_offset_0),
	.prn(vcc));
defparam \ic_fill_ap_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[0] .power_up = "low";

dffeas \ic_fill_line[1] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_1),
	.prn(vcc));
defparam \ic_fill_line[1] .is_wysiwyg = "true";
defparam \ic_fill_line[1] .power_up = "low";

dffeas \ic_fill_line[0] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_0),
	.prn(vcc));
defparam \ic_fill_line[0] .is_wysiwyg = "true";
defparam \ic_fill_line[0] .power_up = "low";

dffeas \ic_fill_ap_offset[2] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[1]~0_combout ),
	.q(ic_fill_ap_offset_2),
	.prn(vcc));
defparam \ic_fill_ap_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[2] .power_up = "low";

dffeas \ic_fill_ap_offset[1] (
	.clk(clk_clk),
	.d(\ic_fill_ap_offset_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[1]~0_combout ),
	.q(ic_fill_ap_offset_1),
	.prn(vcc));
defparam \ic_fill_ap_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_ap_offset[1] .power_up = "low";

dffeas \ic_fill_line[4] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_4),
	.prn(vcc));
defparam \ic_fill_line[4] .is_wysiwyg = "true";
defparam \ic_fill_line[4] .power_up = "low";

dffeas \ic_fill_line[3] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_3),
	.prn(vcc));
defparam \ic_fill_line[3] .is_wysiwyg = "true";
defparam \ic_fill_line[3] .power_up = "low";

dffeas \ic_fill_line[2] (
	.clk(clk_clk),
	.d(\ic_tag_wraddress_nxt~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ic_fill_line_2),
	.prn(vcc));
defparam \ic_fill_line[2] .is_wysiwyg = "true";
defparam \ic_fill_line[2] .power_up = "low";

dffeas \d_byteenable[2]~reg0 (
	.clk(clk_clk),
	.d(\d_byteenable_nxt[2]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_2),
	.prn(vcc));
defparam \d_byteenable[2]~reg0 .is_wysiwyg = "true";
defparam \d_byteenable[2]~reg0 .power_up = "low";

dffeas \d_byteenable[3]~reg0 (
	.clk(clk_clk),
	.d(\d_byteenable_nxt[3]~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(d_byteenable_3),
	.prn(vcc));
defparam \d_byteenable[3]~reg0 .is_wysiwyg = "true";
defparam \d_byteenable[3]~reg0 .power_up = "low";

dffeas \d_writedata[31]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[31]~28_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_31),
	.prn(vcc));
defparam \d_writedata[31]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[31]~reg0 .power_up = "low";

dffeas \d_writedata[29]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[29]~29_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_29),
	.prn(vcc));
defparam \d_writedata[29]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[29]~reg0 .power_up = "low";

dffeas \d_writedata[28]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[28]~30_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_28),
	.prn(vcc));
defparam \d_writedata[28]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[28]~reg0 .power_up = "low";

dffeas \d_writedata[30]~reg0 (
	.clk(clk_clk),
	.d(\d_writedata_nxt[30]~31_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\d_writedata[14]~0_combout ),
	.q(d_writedata_30),
	.prn(vcc));
defparam \d_writedata[30]~reg0 .is_wysiwyg = "true";
defparam \d_writedata[30]~reg0 .power_up = "low";

cyclonev_lcell_comb A_dc_wb_wr_starting(
	.dataa(!d_read),
	.datab(!\A_dc_wb_rd_data_first~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_wr_starting~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_wb_wr_starting.extended_lut = "off";
defparam A_dc_wb_wr_starting.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam A_dc_wb_wr_starting.shared_arith = "off";

cyclonev_lcell_comb \av_wr_data_transfer~0 (
	.dataa(!hold_waitrequest),
	.datab(!d_write),
	.datac(!suppress_change_dest_id),
	.datad(!WideOr0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\av_wr_data_transfer~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \av_wr_data_transfer~0 .extended_lut = "off";
defparam \av_wr_data_transfer~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \av_wr_data_transfer~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_wr_data_cnt_nxt[0]~3 (
	.dataa(!\A_dc_wb_wr_starting~combout ),
	.datab(!\av_wr_data_transfer~0_combout ),
	.datac(!\A_dc_wr_data_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wr_data_cnt_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wr_data_cnt_nxt[0]~3 .extended_lut = "off";
defparam \A_dc_wr_data_cnt_nxt[0]~3 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \A_dc_wr_data_cnt_nxt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \hq3myc14108phmpo7y7qmhbp98hy0vq~0 (
	.dataa(!r_sync_rst),
	.datab(!NJQG9082),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hq3myc14108phmpo7y7qmhbp98hy0vq~0 .extended_lut = "off";
defparam \hq3myc14108phmpo7y7qmhbp98hy0vq~0 .lut_mask = 64'h7777777777777777;
defparam \hq3myc14108phmpo7y7qmhbp98hy0vq~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_wb_wr_active_nxt~0 (
	.dataa(!\A_dc_wb_wr_starting~combout ),
	.datab(!\A_dc_wb_wr_active~q ),
	.datac(!\A_dc_wr_data_cnt[3]~q ),
	.datad(!\av_wr_data_transfer~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_wr_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_wr_active_nxt~0 .extended_lut = "off";
defparam \A_dc_wb_wr_active_nxt~0 .lut_mask = 64'hF7D5F7D5F7D5F7D5;
defparam \A_dc_wb_wr_active_nxt~0 .shared_arith = "off";

dffeas A_dc_wb_wr_active(
	.clk(clk_clk),
	.d(\A_dc_wb_wr_active_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_wb_wr_active~q ),
	.prn(vcc));
defparam A_dc_wb_wr_active.is_wysiwyg = "true";
defparam A_dc_wb_wr_active.power_up = "low";

cyclonev_lcell_comb \A_dc_wr_data_cnt[2]~0 (
	.dataa(!hold_waitrequest),
	.datab(!d_write),
	.datac(!\A_dc_wb_wr_starting~combout ),
	.datad(!\A_dc_wb_wr_active~q ),
	.datae(!suppress_change_dest_id),
	.dataf(!WideOr0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wr_data_cnt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wr_data_cnt[2]~0 .extended_lut = "off";
defparam \A_dc_wr_data_cnt[2]~0 .lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam \A_dc_wr_data_cnt[2]~0 .shared_arith = "off";

dffeas \A_dc_wr_data_cnt[0] (
	.clk(clk_clk),
	.d(\A_dc_wr_data_cnt_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wr_data_cnt[2]~0_combout ),
	.q(\A_dc_wr_data_cnt[0]~q ),
	.prn(vcc));
defparam \A_dc_wr_data_cnt[0] .is_wysiwyg = "true";
defparam \A_dc_wr_data_cnt[0] .power_up = "low";

cyclonev_lcell_comb \A_dc_wr_data_cnt_nxt[1]~2 (
	.dataa(!\av_wr_data_transfer~0_combout ),
	.datab(!\A_dc_wr_data_cnt[1]~q ),
	.datac(!\A_dc_wr_data_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wr_data_cnt_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wr_data_cnt_nxt[1]~2 .extended_lut = "off";
defparam \A_dc_wr_data_cnt_nxt[1]~2 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \A_dc_wr_data_cnt_nxt[1]~2 .shared_arith = "off";

dffeas \A_dc_wr_data_cnt[1] (
	.clk(clk_clk),
	.d(\A_dc_wr_data_cnt_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wr_data_cnt[2]~0_combout ),
	.q(\A_dc_wr_data_cnt[1]~q ),
	.prn(vcc));
defparam \A_dc_wr_data_cnt[1] .is_wysiwyg = "true";
defparam \A_dc_wr_data_cnt[1] .power_up = "low";

cyclonev_lcell_comb \A_dc_wr_data_cnt_nxt[2]~1 (
	.dataa(!\av_wr_data_transfer~0_combout ),
	.datab(!\A_dc_wr_data_cnt[2]~q ),
	.datac(!\A_dc_wr_data_cnt[1]~q ),
	.datad(!\A_dc_wr_data_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wr_data_cnt_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wr_data_cnt_nxt[2]~1 .extended_lut = "off";
defparam \A_dc_wr_data_cnt_nxt[2]~1 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \A_dc_wr_data_cnt_nxt[2]~1 .shared_arith = "off";

dffeas \A_dc_wr_data_cnt[2] (
	.clk(clk_clk),
	.d(\A_dc_wr_data_cnt_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wr_data_cnt[2]~0_combout ),
	.q(\A_dc_wr_data_cnt[2]~q ),
	.prn(vcc));
defparam \A_dc_wr_data_cnt[2] .is_wysiwyg = "true";
defparam \A_dc_wr_data_cnt[2] .power_up = "low";

cyclonev_lcell_comb \A_dc_wr_data_cnt_nxt[3]~0 (
	.dataa(!\A_dc_wb_wr_starting~combout ),
	.datab(!\A_dc_wr_data_cnt[3]~q ),
	.datac(!\av_wr_data_transfer~0_combout ),
	.datad(!\A_dc_wr_data_cnt[2]~q ),
	.datae(!\A_dc_wr_data_cnt[1]~q ),
	.dataf(!\A_dc_wr_data_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wr_data_cnt_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wr_data_cnt_nxt[3]~0 .extended_lut = "off";
defparam \A_dc_wr_data_cnt_nxt[3]~0 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \A_dc_wr_data_cnt_nxt[3]~0 .shared_arith = "off";

dffeas \A_dc_wr_data_cnt[3] (
	.clk(clk_clk),
	.d(\A_dc_wr_data_cnt_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_wr_data_cnt[2]~0_combout ),
	.q(\A_dc_wr_data_cnt[3]~q ),
	.prn(vcc));
defparam \A_dc_wr_data_cnt[3] .is_wysiwyg = "true";
defparam \A_dc_wr_data_cnt[3] .power_up = "low";

cyclonev_lcell_comb \A_dc_wb_active_nxt~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_wr_data_cnt[3]~q ),
	.datac(!\av_wr_data_transfer~0_combout ),
	.datad(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_active_nxt~0 .extended_lut = "off";
defparam \A_dc_wb_active_nxt~0 .lut_mask = 64'hD8FFD8FFD8FFD8FF;
defparam \A_dc_wb_active_nxt~0 .shared_arith = "off";

dffeas A_dc_wb_active(
	.clk(clk_clk),
	.d(\A_dc_wb_active_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_wb_active~q ),
	.prn(vcc));
defparam A_dc_wb_active.is_wysiwyg = "true";
defparam A_dc_wb_active.power_up = "low";

dffeas \E_iw[0] (
	.clk(clk_clk),
	.d(\D_iw[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[0]~q ),
	.prn(vcc));
defparam \E_iw[0] .is_wysiwyg = "true";
defparam \E_iw[0] .power_up = "low";

cyclonev_lcell_comb \F_iw[5]~1 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[5]~1 .extended_lut = "off";
defparam \F_iw[5]~1 .lut_mask = 64'h7777777777777777;
defparam \F_iw[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[3]~2 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[3]~2 .extended_lut = "off";
defparam \F_iw[3]~2 .lut_mask = 64'h7777777777777777;
defparam \F_iw[3]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[1]~3 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[1]~3 .extended_lut = "off";
defparam \F_iw[1]~3 .lut_mask = 64'h7777777777777777;
defparam \F_iw[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[4]~4 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[4]~4 .extended_lut = "off";
defparam \F_iw[4]~4 .lut_mask = 64'h7777777777777777;
defparam \F_iw[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[2]~5 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[2]~5 .extended_lut = "off";
defparam \F_iw[2]~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_a_not_src~0 (
	.dataa(!\F_iw[5]~1_combout ),
	.datab(!\F_iw[3]~2_combout ),
	.datac(!\F_iw[1]~3_combout ),
	.datad(!\F_iw[4]~4_combout ),
	.datae(!\F_iw[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_a_not_src~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_a_not_src~0 .extended_lut = "off";
defparam \F_ctrl_a_not_src~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \F_ctrl_a_not_src~0 .shared_arith = "off";

dffeas D_ctrl_a_not_src(
	.clk(clk_clk),
	.d(\F_ctrl_a_not_src~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_a_not_src~q ),
	.prn(vcc));
defparam D_ctrl_a_not_src.is_wysiwyg = "true";
defparam D_ctrl_a_not_src.power_up = "low";

cyclonev_lcell_comb \F_ctrl_b_is_dst~0 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_b_is_dst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_b_is_dst~0 .extended_lut = "off";
defparam \F_ctrl_b_is_dst~0 .lut_mask = 64'hFFBEFFBEFFBEFFBE;
defparam \F_ctrl_b_is_dst~0 .shared_arith = "off";

dffeas D_ctrl_b_is_dst(
	.clk(clk_clk),
	.d(\F_ctrl_b_is_dst~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_b_is_dst~q ),
	.prn(vcc));
defparam D_ctrl_b_is_dst.is_wysiwyg = "true";
defparam D_ctrl_b_is_dst.power_up = "low";

dffeas M_ctrl_late_result(
	.clk(clk_clk),
	.d(\E_ctrl_late_result~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_late_result~q ),
	.prn(vcc));
defparam M_ctrl_late_result.is_wysiwyg = "true";
defparam M_ctrl_late_result.power_up = "low";

cyclonev_lcell_comb \F_iw[19]~13 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[19] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[19]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[19]~13 .extended_lut = "off";
defparam \F_iw[19]~13 .lut_mask = 64'h7777777777777777;
defparam \F_iw[19]~13 .shared_arith = "off";

dffeas \D_iw[19] (
	.clk(clk_clk),
	.d(\F_iw[19]~13_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[19]~q ),
	.prn(vcc));
defparam \D_iw[19] .is_wysiwyg = "true";
defparam \D_iw[19] .power_up = "low";

dffeas \D_iw[24] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[24]~q ),
	.prn(vcc));
defparam \D_iw[24] .is_wysiwyg = "true";
defparam \D_iw[24] .power_up = "low";

cyclonev_lcell_comb \F_ctrl_implicit_dst_retaddr~0 (
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[5]~1_combout ),
	.datac(!\F_iw[3]~2_combout ),
	.datad(!\F_iw[4]~4_combout ),
	.datae(!\F_iw[2]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_implicit_dst_retaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_implicit_dst_retaddr~0 .extended_lut = "off";
defparam \F_ctrl_implicit_dst_retaddr~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \F_ctrl_implicit_dst_retaddr~0 .shared_arith = "off";

dffeas D_ctrl_implicit_dst_retaddr(
	.clk(clk_clk),
	.d(\F_ctrl_implicit_dst_retaddr~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_implicit_dst_retaddr~q ),
	.prn(vcc));
defparam D_ctrl_implicit_dst_retaddr.is_wysiwyg = "true";
defparam D_ctrl_implicit_dst_retaddr.power_up = "low";

cyclonev_lcell_comb \F_iw[13]~8 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[13]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[13]~8 .extended_lut = "off";
defparam \F_iw[13]~8 .lut_mask = 64'h7777777777777777;
defparam \F_iw[13]~8 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_implicit_dst_eretaddr~0 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.datac(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datae(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_implicit_dst_eretaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_implicit_dst_eretaddr~0 .extended_lut = "off";
defparam \F_ctrl_implicit_dst_eretaddr~0 .lut_mask = 64'hFEFFEFFFEFFFFEFF;
defparam \F_ctrl_implicit_dst_eretaddr~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal2~0 (
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[5]~1_combout ),
	.datac(!\F_iw[3]~2_combout ),
	.datad(!\F_iw[1]~3_combout ),
	.datae(!\F_iw[4]~4_combout ),
	.dataf(!\F_iw[2]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal2~0 .extended_lut = "off";
defparam \Equal2~0 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \Equal2~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_implicit_dst_eretaddr~1 (
	.dataa(!\F_iw[13]~8_combout ),
	.datab(!\F_ctrl_implicit_dst_eretaddr~0_combout ),
	.datac(!\Equal2~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_implicit_dst_eretaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_implicit_dst_eretaddr~1 .extended_lut = "off";
defparam \F_ctrl_implicit_dst_eretaddr~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \F_ctrl_implicit_dst_eretaddr~1 .shared_arith = "off";

dffeas D_ctrl_implicit_dst_eretaddr(
	.clk(clk_clk),
	.d(\F_ctrl_implicit_dst_eretaddr~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_implicit_dst_eretaddr~q ),
	.prn(vcc));
defparam D_ctrl_implicit_dst_eretaddr.is_wysiwyg = "true";
defparam D_ctrl_implicit_dst_eretaddr.power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[2]~3 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[19]~q ),
	.datac(!\D_iw[24]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[2]~3 .extended_lut = "off";
defparam \D_dst_regnum[2]~3 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[2]~3 .shared_arith = "off";

dffeas \E_dst_regnum[2] (
	.clk(clk_clk),
	.d(\D_dst_regnum[2]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_dst_regnum[2]~q ),
	.prn(vcc));
defparam \E_dst_regnum[2] .is_wysiwyg = "true";
defparam \E_dst_regnum[2] .power_up = "low";

cyclonev_lcell_comb \F_iw[16]~6 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[16]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[16]~6 .extended_lut = "off";
defparam \F_iw[16]~6 .lut_mask = 64'h7777777777777777;
defparam \F_iw[16]~6 .shared_arith = "off";

dffeas \D_iw[16] (
	.clk(clk_clk),
	.d(\F_iw[16]~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[16]~q ),
	.prn(vcc));
defparam \D_iw[16] .is_wysiwyg = "true";
defparam \D_iw[16] .power_up = "low";

dffeas \E_iw[16] (
	.clk(clk_clk),
	.d(\D_iw[16]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[16]~q ),
	.prn(vcc));
defparam \E_iw[16] .is_wysiwyg = "true";
defparam \E_iw[16] .power_up = "low";

cyclonev_lcell_comb \F_iw[15]~7 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[15]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[15]~7 .extended_lut = "off";
defparam \F_iw[15]~7 .lut_mask = 64'h7777777777777777;
defparam \F_iw[15]~7 .shared_arith = "off";

dffeas \D_iw[15] (
	.clk(clk_clk),
	.d(\F_iw[15]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[15]~q ),
	.prn(vcc));
defparam \D_iw[15] .is_wysiwyg = "true";
defparam \D_iw[15] .power_up = "low";

dffeas \E_iw[15] (
	.clk(clk_clk),
	.d(\D_iw[15]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[15]~q ),
	.prn(vcc));
defparam \E_iw[15] .is_wysiwyg = "true";
defparam \E_iw[15] .power_up = "low";

dffeas \D_iw[13] (
	.clk(clk_clk),
	.d(\F_iw[13]~8_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[13]~q ),
	.prn(vcc));
defparam \D_iw[13] .is_wysiwyg = "true";
defparam \D_iw[13] .power_up = "low";

dffeas \E_iw[13] (
	.clk(clk_clk),
	.d(\D_iw[13]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[13]~q ),
	.prn(vcc));
defparam \E_iw[13] .is_wysiwyg = "true";
defparam \E_iw[13] .power_up = "low";

cyclonev_lcell_comb \E_hbreak_req~0 (
	.dataa(!\E_iw[16]~q ),
	.datab(!\E_iw[15]~q ),
	.datac(!\E_iw[13]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_hbreak_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_hbreak_req~0 .extended_lut = "off";
defparam \E_hbreak_req~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_hbreak_req~0 .shared_arith = "off";

dffeas \D_iw[3] (
	.clk(clk_clk),
	.d(\F_iw[3]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[3]~q ),
	.prn(vcc));
defparam \D_iw[3] .is_wysiwyg = "true";
defparam \D_iw[3] .power_up = "low";

dffeas \E_iw[3] (
	.clk(clk_clk),
	.d(\D_iw[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[3]~q ),
	.prn(vcc));
defparam \E_iw[3] .is_wysiwyg = "true";
defparam \E_iw[3] .power_up = "low";

dffeas \D_iw[1] (
	.clk(clk_clk),
	.d(\F_iw[1]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[1]~q ),
	.prn(vcc));
defparam \D_iw[1] .is_wysiwyg = "true";
defparam \D_iw[1] .power_up = "low";

dffeas \E_iw[1] (
	.clk(clk_clk),
	.d(\D_iw[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[1]~q ),
	.prn(vcc));
defparam \E_iw[1] .is_wysiwyg = "true";
defparam \E_iw[1] .power_up = "low";

dffeas \D_iw[4] (
	.clk(clk_clk),
	.d(\F_iw[4]~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[4]~q ),
	.prn(vcc));
defparam \D_iw[4] .is_wysiwyg = "true";
defparam \D_iw[4] .power_up = "low";

dffeas \E_iw[4] (
	.clk(clk_clk),
	.d(\D_iw[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[4]~q ),
	.prn(vcc));
defparam \E_iw[4] .is_wysiwyg = "true";
defparam \E_iw[4] .power_up = "low";

dffeas \D_iw[2] (
	.clk(clk_clk),
	.d(\F_iw[2]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[2]~q ),
	.prn(vcc));
defparam \D_iw[2] .is_wysiwyg = "true";
defparam \D_iw[2] .power_up = "low";

dffeas \E_iw[2] (
	.clk(clk_clk),
	.d(\D_iw[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[2]~q ),
	.prn(vcc));
defparam \E_iw[2] .is_wysiwyg = "true";
defparam \E_iw[2] .power_up = "low";

cyclonev_lcell_comb \Equal209~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[3]~q ),
	.datad(!\E_iw[1]~q ),
	.datae(!\E_iw[4]~q ),
	.dataf(!\E_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal209~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal209~0 .extended_lut = "off";
defparam \Equal209~0 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \Equal209~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[14]~10 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[14]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[14]~10 .extended_lut = "off";
defparam \F_iw[14]~10 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[14]~10 .shared_arith = "off";

dffeas \D_iw[14] (
	.clk(clk_clk),
	.d(\F_iw[14]~10_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[14]~q ),
	.prn(vcc));
defparam \D_iw[14] .is_wysiwyg = "true";
defparam \D_iw[14] .power_up = "low";

dffeas \E_iw[14] (
	.clk(clk_clk),
	.d(\D_iw[14]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[14]~q ),
	.prn(vcc));
defparam \E_iw[14] .is_wysiwyg = "true";
defparam \E_iw[14] .power_up = "low";

cyclonev_lcell_comb \F_iw[12]~11 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[12]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[12]~11 .extended_lut = "off";
defparam \F_iw[12]~11 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[12]~11 .shared_arith = "off";

dffeas \D_iw[12] (
	.clk(clk_clk),
	.d(\F_iw[12]~11_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[12]~q ),
	.prn(vcc));
defparam \D_iw[12] .is_wysiwyg = "true";
defparam \D_iw[12] .power_up = "low";

dffeas \E_iw[12] (
	.clk(clk_clk),
	.d(\D_iw[12]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[12]~q ),
	.prn(vcc));
defparam \E_iw[12] .is_wysiwyg = "true";
defparam \E_iw[12] .power_up = "low";

cyclonev_lcell_comb \F_iw[11]~12 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[11]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[11]~12 .extended_lut = "off";
defparam \F_iw[11]~12 .lut_mask = 64'h7777777777777777;
defparam \F_iw[11]~12 .shared_arith = "off";

dffeas \D_iw[11] (
	.clk(clk_clk),
	.d(\F_iw[11]~12_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[11]~q ),
	.prn(vcc));
defparam \D_iw[11] .is_wysiwyg = "true";
defparam \D_iw[11] .power_up = "low";

dffeas \E_iw[11] (
	.clk(clk_clk),
	.d(\D_iw[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[11]~q ),
	.prn(vcc));
defparam \E_iw[11] .is_wysiwyg = "true";
defparam \E_iw[11] .power_up = "low";

cyclonev_lcell_comb \E_hbreak_req~1 (
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_iw[12]~q ),
	.datac(!\E_iw[11]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_hbreak_req~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_hbreak_req~1 .extended_lut = "off";
defparam \E_hbreak_req~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \E_hbreak_req~1 .shared_arith = "off";

cyclonev_lcell_comb E_hbreak_req(
	.dataa(!\E_valid~0_combout ),
	.datab(!\E_hbreak_req~0_combout ),
	.datac(!\Equal209~0_combout ),
	.datad(!\E_hbreak_req~1_combout ),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_hbreak_req~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_hbreak_req.extended_lut = "off";
defparam E_hbreak_req.lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam E_hbreak_req.shared_arith = "off";

dffeas \D_bht_data[1] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_bht|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_bht_data[1]~q ),
	.prn(vcc));
defparam \D_bht_data[1] .is_wysiwyg = "true";
defparam \D_bht_data[1] .power_up = "low";

dffeas \E_bht_data[1] (
	.clk(clk_clk),
	.d(\D_bht_data[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_bht_data[1]~q ),
	.prn(vcc));
defparam \E_bht_data[1] .is_wysiwyg = "true";
defparam \E_bht_data[1] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_cmp~3 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[12]~q ),
	.datae(!\D_iw[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~3 .extended_lut = "off";
defparam \D_ctrl_cmp~3 .lut_mask = 64'hFFFFFFF6FFFFFFF6;
defparam \D_ctrl_cmp~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[15]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~0 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \D_ctrl_alu_subtract~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~1 (
	.dataa(!\D_iw[0]~q ),
	.datab(gnd),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~1 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~1 .lut_mask = 64'hAFFAFAAFFAAFAFFA;
defparam \D_ctrl_alu_subtract~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_subtract~2 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\Equal171~0_combout ),
	.datac(!\D_ctrl_cmp~3_combout ),
	.datad(!\D_ctrl_alu_subtract~0_combout ),
	.datae(!\D_ctrl_alu_subtract~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_subtract~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_subtract~2 .extended_lut = "off";
defparam \D_ctrl_alu_subtract~2 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \D_ctrl_alu_subtract~2 .shared_arith = "off";

dffeas E_ctrl_alu_subtract(
	.clk(clk_clk),
	.d(\D_ctrl_alu_subtract~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_alu_subtract~q ),
	.prn(vcc));
defparam E_ctrl_alu_subtract.is_wysiwyg = "true";
defparam E_ctrl_alu_subtract.power_up = "low";

cyclonev_lcell_comb \Equal154~1 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal154~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal154~1 .extended_lut = "off";
defparam \Equal154~1 .lut_mask = 64'hFFFFFFFFFFFFFEFF;
defparam \Equal154~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal154~3 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal154~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal154~3 .extended_lut = "off";
defparam \Equal154~3 .lut_mask = 64'hFFFFFFFFFFFEFFFF;
defparam \Equal154~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_signed_comparison~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_signed_comparison~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_signed_comparison~0 .extended_lut = "off";
defparam \D_ctrl_alu_signed_comparison~0 .lut_mask = 64'hEFFEFEEFFEEFEFFE;
defparam \D_ctrl_alu_signed_comparison~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_signed_comparison~1 (
	.dataa(!\Equal171~0_combout ),
	.datab(!\Equal154~1_combout ),
	.datac(!\Equal154~3_combout ),
	.datad(!\D_ctrl_alu_signed_comparison~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_signed_comparison~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_signed_comparison~1 .extended_lut = "off";
defparam \D_ctrl_alu_signed_comparison~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_alu_signed_comparison~1 .shared_arith = "off";

dffeas E_ctrl_alu_signed_comparison(
	.clk(clk_clk),
	.d(\D_ctrl_alu_signed_comparison~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_alu_signed_comparison~q ),
	.prn(vcc));
defparam E_ctrl_alu_signed_comparison.is_wysiwyg = "true";
defparam E_ctrl_alu_signed_comparison.power_up = "low";

cyclonev_lcell_comb \F_ctrl_src2_choose_imm~0 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datac(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_src2_choose_imm~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_src2_choose_imm~0 .extended_lut = "off";
defparam \F_ctrl_src2_choose_imm~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \F_ctrl_src2_choose_imm~0 .shared_arith = "off";

cyclonev_lcell_comb F_ctrl_src2_choose_imm(
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datad(!\F_iw[12]~11_combout ),
	.datae(!\Equal2~0_combout ),
	.dataf(!\F_ctrl_src2_choose_imm~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_src2_choose_imm~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_ctrl_src2_choose_imm.extended_lut = "off";
defparam F_ctrl_src2_choose_imm.lut_mask = 64'hFBFFFFFFFFFFFFFF;
defparam F_ctrl_src2_choose_imm.shared_arith = "off";

dffeas D_ctrl_src2_choose_imm(
	.clk(clk_clk),
	.d(\F_ctrl_src2_choose_imm~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_src2_choose_imm~q ),
	.prn(vcc));
defparam D_ctrl_src2_choose_imm.is_wysiwyg = "true";
defparam D_ctrl_src2_choose_imm.power_up = "low";

dffeas \D_iw[23] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[23]~q ),
	.prn(vcc));
defparam \D_iw[23] .is_wysiwyg = "true";
defparam \D_iw[23] .power_up = "low";

cyclonev_lcell_comb \F_iw[18]~14 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[18] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[18]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[18]~14 .extended_lut = "off";
defparam \F_iw[18]~14 .lut_mask = 64'h7777777777777777;
defparam \F_iw[18]~14 .shared_arith = "off";

dffeas \D_iw[18] (
	.clk(clk_clk),
	.d(\F_iw[18]~14_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[18]~q ),
	.prn(vcc));
defparam \D_iw[18] .is_wysiwyg = "true";
defparam \D_iw[18] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[1]~0 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[23]~q ),
	.datac(!\D_iw[18]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[1]~0 .extended_lut = "off";
defparam \D_dst_regnum[1]~0 .lut_mask = 64'hBFFF1FFFBFFF1FFF;
defparam \D_dst_regnum[1]~0 .shared_arith = "off";

dffeas \D_iw[26] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[26]~q ),
	.prn(vcc));
defparam \D_iw[26] .is_wysiwyg = "true";
defparam \D_iw[26] .power_up = "low";

cyclonev_lcell_comb \F_iw[21]~15 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[21] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[21]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[21]~15 .extended_lut = "off";
defparam \F_iw[21]~15 .lut_mask = 64'h7777777777777777;
defparam \F_iw[21]~15 .shared_arith = "off";

dffeas \D_iw[21] (
	.clk(clk_clk),
	.d(\F_iw[21]~15_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[21]~q ),
	.prn(vcc));
defparam \D_iw[21] .is_wysiwyg = "true";
defparam \D_iw[21] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[4]~1 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[26]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[4]~1 .extended_lut = "off";
defparam \D_dst_regnum[4]~1 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[4]~1 .shared_arith = "off";

cyclonev_lcell_comb F_ctrl_ignore_dst(
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[1]~3_combout ),
	.datac(!\F_iw[2]~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_ignore_dst~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_ctrl_ignore_dst.extended_lut = "off";
defparam F_ctrl_ignore_dst.lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam F_ctrl_ignore_dst.shared_arith = "off";

dffeas D_ctrl_ignore_dst(
	.clk(clk_clk),
	.d(\F_ctrl_ignore_dst~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_ignore_dst~q ),
	.prn(vcc));
defparam D_ctrl_ignore_dst.is_wysiwyg = "true";
defparam D_ctrl_ignore_dst.power_up = "low";

dffeas \D_iw[22] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[22]~q ),
	.prn(vcc));
defparam \D_iw[22] .is_wysiwyg = "true";
defparam \D_iw[22] .power_up = "low";

dffeas \D_iw[17] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[17]~q ),
	.prn(vcc));
defparam \D_iw[17] .is_wysiwyg = "true";
defparam \D_iw[17] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[0]~2 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[22]~q ),
	.datac(!\D_iw[17]~q ),
	.datad(!\D_ctrl_implicit_dst_retaddr~q ),
	.datae(!\D_ctrl_implicit_dst_eretaddr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[0]~2 .extended_lut = "off";
defparam \D_dst_regnum[0]~2 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[0]~2 .shared_arith = "off";

dffeas \D_iw[25] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[25]~q ),
	.prn(vcc));
defparam \D_iw[25] .is_wysiwyg = "true";
defparam \D_iw[25] .power_up = "low";

cyclonev_lcell_comb \F_iw[20]~16 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[20] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[20]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[20]~16 .extended_lut = "off";
defparam \F_iw[20]~16 .lut_mask = 64'h7777777777777777;
defparam \F_iw[20]~16 .shared_arith = "off";

dffeas \D_iw[20] (
	.clk(clk_clk),
	.d(\F_iw[20]~16_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[20]~q ),
	.prn(vcc));
defparam \D_iw[20] .is_wysiwyg = "true";
defparam \D_iw[20] .power_up = "low";

cyclonev_lcell_comb \D_dst_regnum[3]~4 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\D_iw[25]~q ),
	.datac(!\D_ctrl_implicit_dst_retaddr~q ),
	.datad(!\D_ctrl_implicit_dst_eretaddr~q ),
	.datae(!\D_iw[20]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dst_regnum[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dst_regnum[3]~4 .extended_lut = "off";
defparam \D_dst_regnum[3]~4 .lut_mask = 64'h27FFFFFF27FFFFFF;
defparam \D_dst_regnum[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal295~0 (
	.dataa(!\D_dst_regnum[0]~2_combout ),
	.datab(!\D_dst_regnum[2]~3_combout ),
	.datac(!\D_dst_regnum[3]~4_combout ),
	.datad(!\D_dst_regnum[4]~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal295~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal295~0 .extended_lut = "off";
defparam \Equal295~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal295~0 .shared_arith = "off";

cyclonev_lcell_comb D_wr_dst_reg(
	.dataa(!\D_valid~combout ),
	.datab(!\D_ctrl_ignore_dst~q ),
	.datac(!\D_dst_regnum[1]~0_combout ),
	.datad(!\Equal295~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_wr_dst_reg~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_wr_dst_reg.extended_lut = "off";
defparam D_wr_dst_reg.lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam D_wr_dst_reg.shared_arith = "off";

cyclonev_lcell_comb \D_regnum_b_cmp_F~0 (
	.dataa(!\D_dst_regnum[0]~2_combout ),
	.datab(!\D_dst_regnum[2]~3_combout ),
	.datac(!\D_dst_regnum[3]~4_combout ),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datae(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \D_regnum_b_cmp_F~0 .lut_mask = 64'h6996966996696996;
defparam \D_regnum_b_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb D_regnum_b_cmp_F(
	.dataa(!\D_dst_regnum[1]~0_combout ),
	.datab(!\D_dst_regnum[4]~1_combout ),
	.datac(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datae(!\D_wr_dst_reg~combout ),
	.dataf(!\D_regnum_b_cmp_F~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_regnum_b_cmp_F.extended_lut = "off";
defparam D_regnum_b_cmp_F.lut_mask = 64'h6996FFFFFFFFFFFF;
defparam D_regnum_b_cmp_F.shared_arith = "off";

dffeas E_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\D_regnum_b_cmp_F~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_stall~combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam E_regnum_b_cmp_D.is_wysiwyg = "true";
defparam E_regnum_b_cmp_D.power_up = "low";

dffeas \E_dst_regnum[4] (
	.clk(clk_clk),
	.d(\D_dst_regnum[4]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_dst_regnum[4]~q ),
	.prn(vcc));
defparam \E_dst_regnum[4] .is_wysiwyg = "true";
defparam \E_dst_regnum[4] .power_up = "low";

dffeas \M_dst_regnum[4] (
	.clk(clk_clk),
	.d(\E_dst_regnum[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_dst_regnum[4]~q ),
	.prn(vcc));
defparam \M_dst_regnum[4] .is_wysiwyg = "true";
defparam \M_dst_regnum[4] .power_up = "low";

dffeas M_wr_dst_reg_from_E(
	.clk(clk_clk),
	.d(\E_wr_dst_reg~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_wr_dst_reg_from_E~q ),
	.prn(vcc));
defparam M_wr_dst_reg_from_E.is_wysiwyg = "true";
defparam M_wr_dst_reg_from_E.power_up = "low";

dffeas \E_dst_regnum[0] (
	.clk(clk_clk),
	.d(\D_dst_regnum[0]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_dst_regnum[0]~q ),
	.prn(vcc));
defparam \E_dst_regnum[0] .is_wysiwyg = "true";
defparam \E_dst_regnum[0] .power_up = "low";

dffeas \M_dst_regnum[0] (
	.clk(clk_clk),
	.d(\E_dst_regnum[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_dst_regnum[0]~q ),
	.prn(vcc));
defparam \M_dst_regnum[0] .is_wysiwyg = "true";
defparam \M_dst_regnum[0] .power_up = "low";

dffeas \E_dst_regnum[1] (
	.clk(clk_clk),
	.d(\D_dst_regnum[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_dst_regnum[1]~q ),
	.prn(vcc));
defparam \E_dst_regnum[1] .is_wysiwyg = "true";
defparam \E_dst_regnum[1] .power_up = "low";

dffeas \M_dst_regnum[1] (
	.clk(clk_clk),
	.d(\E_dst_regnum[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_dst_regnum[1]~q ),
	.prn(vcc));
defparam \M_dst_regnum[1] .is_wysiwyg = "true";
defparam \M_dst_regnum[1] .power_up = "low";

cyclonev_lcell_comb \M_regnum_b_cmp_F~0 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\M_wr_dst_reg_from_E~q ),
	.datad(!\M_dst_regnum[0]~q ),
	.datae(!\M_dst_regnum[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \M_regnum_b_cmp_F~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \M_regnum_b_cmp_F~0 .shared_arith = "off";

dffeas \M_dst_regnum[2] (
	.clk(clk_clk),
	.d(\E_dst_regnum[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_dst_regnum[2]~q ),
	.prn(vcc));
defparam \M_dst_regnum[2] .is_wysiwyg = "true";
defparam \M_dst_regnum[2] .power_up = "low";

dffeas \E_dst_regnum[3] (
	.clk(clk_clk),
	.d(\D_dst_regnum[3]~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_dst_regnum[3]~q ),
	.prn(vcc));
defparam \E_dst_regnum[3] .is_wysiwyg = "true";
defparam \E_dst_regnum[3] .power_up = "low";

dffeas \M_dst_regnum[3] (
	.clk(clk_clk),
	.d(\E_dst_regnum[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_dst_regnum[3]~q ),
	.prn(vcc));
defparam \M_dst_regnum[3] .is_wysiwyg = "true";
defparam \M_dst_regnum[3] .power_up = "low";

cyclonev_lcell_comb \M_regnum_b_cmp_F~1 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datac(!\M_dst_regnum[2]~q ),
	.datad(!\M_dst_regnum[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_b_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_b_cmp_F~1 .extended_lut = "off";
defparam \M_regnum_b_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \M_regnum_b_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb M_regnum_b_cmp_F(
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datab(!\M_dst_regnum[4]~q ),
	.datac(!\M_regnum_b_cmp_F~0_combout ),
	.datad(!\M_regnum_b_cmp_F~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_regnum_b_cmp_F.extended_lut = "off";
defparam M_regnum_b_cmp_F.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam M_regnum_b_cmp_F.shared_arith = "off";

dffeas A_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\M_regnum_b_cmp_F~combout ),
	.asdata(\M_regnum_b_cmp_D~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(\A_stall~combout ),
	.q(\A_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam A_regnum_b_cmp_D.is_wysiwyg = "true";
defparam A_regnum_b_cmp_D.power_up = "low";

dffeas \A_dst_regnum_from_M[4] (
	.clk(clk_clk),
	.d(\M_dst_regnum[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dst_regnum_from_M[4]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[4] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[4] .power_up = "low";

dffeas A_wr_dst_reg_from_M(
	.clk(clk_clk),
	.d(\M_wr_dst_reg_from_E~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_wr_dst_reg_from_M~q ),
	.prn(vcc));
defparam A_wr_dst_reg_from_M.is_wysiwyg = "true";
defparam A_wr_dst_reg_from_M.power_up = "low";

dffeas \A_dst_regnum_from_M[0] (
	.clk(clk_clk),
	.d(\M_dst_regnum[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dst_regnum_from_M[0]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[0] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[0] .power_up = "low";

dffeas \A_dst_regnum_from_M[1] (
	.clk(clk_clk),
	.d(\M_dst_regnum[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dst_regnum_from_M[1]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[1] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[1] .power_up = "low";

cyclonev_lcell_comb \A_regnum_b_cmp_F~0 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\A_wr_dst_reg_from_M~q ),
	.datad(!\A_dst_regnum_from_M[0]~q ),
	.datae(!\A_dst_regnum_from_M[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \A_regnum_b_cmp_F~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \A_regnum_b_cmp_F~0 .shared_arith = "off";

dffeas \A_dst_regnum_from_M[2] (
	.clk(clk_clk),
	.d(\M_dst_regnum[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dst_regnum_from_M[2]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[2] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[2] .power_up = "low";

dffeas \A_dst_regnum_from_M[3] (
	.clk(clk_clk),
	.d(\M_dst_regnum[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dst_regnum_from_M[3]~q ),
	.prn(vcc));
defparam \A_dst_regnum_from_M[3] .is_wysiwyg = "true";
defparam \A_dst_regnum_from_M[3] .power_up = "low";

cyclonev_lcell_comb \A_regnum_b_cmp_F~1 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datac(!\A_dst_regnum_from_M[2]~q ),
	.datad(!\A_dst_regnum_from_M[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_b_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_b_cmp_F~1 .extended_lut = "off";
defparam \A_regnum_b_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \A_regnum_b_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb A_regnum_b_cmp_F(
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datab(!\A_dst_regnum_from_M[4]~q ),
	.datac(!\A_regnum_b_cmp_F~0_combout ),
	.datad(!\A_regnum_b_cmp_F~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_regnum_b_cmp_F.extended_lut = "off";
defparam A_regnum_b_cmp_F.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam A_regnum_b_cmp_F.shared_arith = "off";

dffeas W_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\A_regnum_b_cmp_F~combout ),
	.asdata(\A_regnum_b_cmp_D~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(vcc),
	.q(\W_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam W_regnum_b_cmp_D.is_wysiwyg = "true";
defparam W_regnum_b_cmp_D.power_up = "low";

cyclonev_lcell_comb \D_src2_reg[5]~0 (
	.dataa(!\M_regnum_b_cmp_D~q ),
	.datab(!\A_regnum_b_cmp_D~q ),
	.datac(!\W_regnum_b_cmp_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~0 .extended_lut = "off";
defparam \D_src2_reg[5]~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \D_src2_reg[5]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal297~0 (
	.dataa(!\D_iw[26]~q ),
	.datab(!\D_iw[22]~q ),
	.datac(!\D_iw[23]~q ),
	.datad(!\D_iw[24]~q ),
	.datae(!\D_iw[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal297~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal297~0 .extended_lut = "off";
defparam \Equal297~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal297~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[5]~1 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~1 .extended_lut = "off";
defparam \D_src2_reg[5]~1 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \D_src2_reg[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[5]~2 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~2 .extended_lut = "off";
defparam \D_src2_reg[5]~2 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \D_src2_reg[5]~2 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~55 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~55 .extended_lut = "off";
defparam \D_src2_reg[0]~55 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \D_src2_reg[0]~55 .shared_arith = "off";

cyclonev_lcell_comb \Equal92~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[1]~q ),
	.datac(!\D_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal92~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal92~0 .extended_lut = "off";
defparam \Equal92~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \Equal92~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~0 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\Equal171~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~0 .extended_lut = "off";
defparam \D_ctrl_logic~0 .lut_mask = 64'h7777777777777777;
defparam \D_ctrl_logic~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~1 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[11]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_ctrl_logic~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~1 .extended_lut = "off";
defparam \D_ctrl_logic~1 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \D_ctrl_logic~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_logic~2 (
	.dataa(!\D_iw[3]~q ),
	.datab(!\D_iw[4]~q ),
	.datac(!\Equal92~0_combout ),
	.datad(!\D_ctrl_logic~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_logic~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_logic~2 .extended_lut = "off";
defparam \D_ctrl_logic~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_logic~2 .shared_arith = "off";

dffeas E_ctrl_logic(
	.clk(clk_clk),
	.d(\D_ctrl_logic~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_logic~q ),
	.prn(vcc));
defparam E_ctrl_logic.is_wysiwyg = "true";
defparam E_ctrl_logic.power_up = "low";

cyclonev_lcell_comb \Equal105~0 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\D_iw[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal105~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal105~0 .extended_lut = "off";
defparam \Equal105~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \Equal105~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal154~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal154~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal154~0 .extended_lut = "off";
defparam \Equal154~0 .lut_mask = 64'hDFFFFFFFFFFFFFFF;
defparam \Equal154~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~1 .extended_lut = "off";
defparam \D_ctrl_retaddr~1 .lut_mask = 64'h96FF69FF69FF96FF;
defparam \D_ctrl_retaddr~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_retaddr~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\Equal171~0_combout ),
	.datac(!\Equal105~0_combout ),
	.datad(!\Equal154~0_combout ),
	.datae(!\D_ctrl_retaddr~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_retaddr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_retaddr~0 .extended_lut = "off";
defparam \D_ctrl_retaddr~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \D_ctrl_retaddr~0 .shared_arith = "off";

dffeas E_ctrl_retaddr(
	.clk(clk_clk),
	.d(\D_ctrl_retaddr~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_retaddr~q ),
	.prn(vcc));
defparam E_ctrl_retaddr.is_wysiwyg = "true";
defparam E_ctrl_retaddr.power_up = "low";

cyclonev_lcell_comb \D_ctrl_cmp~2 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_iw[14]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[12]~q ),
	.datae(!\D_iw[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~2 .extended_lut = "off";
defparam \D_ctrl_cmp~2 .lut_mask = 64'hFFFFFFF6FFFFFFF6;
defparam \D_ctrl_cmp~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~0 .extended_lut = "off";
defparam \D_ctrl_cmp~0 .lut_mask = 64'hFFFFFFFFFFEBFFBE;
defparam \D_ctrl_cmp~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_cmp~1 (
	.dataa(!\Equal171~0_combout ),
	.datab(!\D_ctrl_cmp~3_combout ),
	.datac(!\D_ctrl_cmp~2_combout ),
	.datad(!\D_ctrl_cmp~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_cmp~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_cmp~1 .extended_lut = "off";
defparam \D_ctrl_cmp~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_cmp~1 .shared_arith = "off";

dffeas E_ctrl_cmp(
	.clk(clk_clk),
	.d(\D_ctrl_cmp~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_cmp~q ),
	.prn(vcc));
defparam E_ctrl_cmp.is_wysiwyg = "true";
defparam E_ctrl_cmp.power_up = "low";

cyclonev_lcell_comb \E_alu_result~0 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_ctrl_cmp~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~0 .extended_lut = "off";
defparam \E_alu_result~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_alu_result~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~3 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(!\D_iw[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~3 .extended_lut = "off";
defparam \D_ctrl_late_result~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_late_result~3 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_mul_lsw~0 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[4]~q ),
	.datad(!\Equal171~0_combout ),
	.datae(!\Equal92~0_combout ),
	.dataf(!\D_ctrl_late_result~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_mul_lsw~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_mul_lsw~0 .extended_lut = "off";
defparam \D_ctrl_mul_lsw~0 .lut_mask = 64'hFDFFFFFFFFFFFFFF;
defparam \D_ctrl_mul_lsw~0 .shared_arith = "off";

dffeas E_ctrl_mul_lsw(
	.clk(clk_clk),
	.d(\D_ctrl_mul_lsw~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_mul_lsw~q ),
	.prn(vcc));
defparam E_ctrl_mul_lsw.is_wysiwyg = "true";
defparam E_ctrl_mul_lsw.power_up = "low";

dffeas M_ctrl_mul_lsw(
	.clk(clk_clk),
	.d(\E_ctrl_mul_lsw~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_mul_lsw~q ),
	.prn(vcc));
defparam M_ctrl_mul_lsw.is_wysiwyg = "true";
defparam M_ctrl_mul_lsw.power_up = "low";

dffeas A_ctrl_mul_lsw(
	.clk(clk_clk),
	.d(\M_ctrl_mul_lsw~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_mul_lsw~q ),
	.prn(vcc));
defparam A_ctrl_mul_lsw.is_wysiwyg = "true";
defparam A_ctrl_mul_lsw.power_up = "low";

cyclonev_lcell_comb \D_logic_op_raw[1]~0 (
	.dataa(!\D_iw[4]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\Equal171~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op_raw[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op_raw[1]~0 .extended_lut = "off";
defparam \D_logic_op_raw[1]~0 .lut_mask = 64'h5353535353535353;
defparam \D_logic_op_raw[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal154~2 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal154~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal154~2 .extended_lut = "off";
defparam \Equal154~2 .lut_mask = 64'hFFFFFEFFFFFFFFFF;
defparam \Equal154~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal154~4 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal154~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal154~4 .extended_lut = "off";
defparam \Equal154~4 .lut_mask = 64'hFFFFFFFFFEFFFFFF;
defparam \Equal154~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal154~5 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal154~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal154~5 .extended_lut = "off";
defparam \Equal154~5 .lut_mask = 64'hFFFFFFFEFFFFFFFF;
defparam \Equal154~5 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~0 (
	.dataa(!\Equal154~1_combout ),
	.datab(!\Equal154~2_combout ),
	.datac(!\Equal154~4_combout ),
	.datad(!\Equal154~5_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~0 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_ctrl_alu_force_xor~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~1 (
	.dataa(!\D_iw[5]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\D_iw[1]~q ),
	.datad(!\D_iw[4]~q ),
	.datae(!\D_iw[2]~q ),
	.dataf(!\D_ctrl_alu_force_xor~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~1 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~1 .lut_mask = 64'hFFFFFFFFFFB7FF7B;
defparam \D_ctrl_alu_force_xor~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_alu_force_xor~2 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_ctrl_alu_force_xor~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_alu_force_xor~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_alu_force_xor~2 .extended_lut = "off";
defparam \D_ctrl_alu_force_xor~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \D_ctrl_alu_force_xor~2 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op[1]~0 (
	.dataa(!\D_logic_op_raw[1]~0_combout ),
	.datab(!\D_ctrl_alu_force_xor~2_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op[1]~0 .extended_lut = "off";
defparam \D_logic_op[1]~0 .lut_mask = 64'h7777777777777777;
defparam \D_logic_op[1]~0 .shared_arith = "off";

dffeas \E_logic_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_logic_op[1]~q ),
	.prn(vcc));
defparam \E_logic_op[1] .is_wysiwyg = "true";
defparam \E_logic_op[1] .power_up = "low";

cyclonev_lcell_comb \D_logic_op_raw[0]~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[3]~q ),
	.datac(!\Equal171~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op_raw[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op_raw[0]~1 .extended_lut = "off";
defparam \D_logic_op_raw[0]~1 .lut_mask = 64'h5353535353535353;
defparam \D_logic_op_raw[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_logic_op[0]~1 (
	.dataa(!\D_ctrl_alu_force_xor~2_combout ),
	.datab(!\D_logic_op_raw[0]~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_logic_op[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_logic_op[0]~1 .extended_lut = "off";
defparam \D_logic_op[0]~1 .lut_mask = 64'h7777777777777777;
defparam \D_logic_op[0]~1 .shared_arith = "off";

dffeas \E_logic_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op[0]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_logic_op[0]~q ),
	.prn(vcc));
defparam \E_logic_op[0] .is_wysiwyg = "true";
defparam \E_logic_op[0] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[31]~9 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[31]~q ),
	.datad(!\E_src1[31]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[31]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[31]~9 .extended_lut = "off";
defparam \E_logic_result[31]~9 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[31]~9 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~30 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[31]~9_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~30 .extended_lut = "off";
defparam \E_alu_result~30 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~30 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[31] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add17~37_sumout ),
	.datac(!\E_alu_result~30_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[31]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[31] .extended_lut = "off";
defparam \E_alu_result[31] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[31] .shared_arith = "off";

dffeas \M_alu_result[31] (
	.clk(clk_clk),
	.d(\E_alu_result[31]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[31]~q ),
	.prn(vcc));
defparam \M_alu_result[31] .is_wysiwyg = "true";
defparam \M_alu_result[31] .power_up = "low";

cyclonev_lcell_comb \E_op_rdctl~0 (
	.dataa(!\E_iw[12]~q ),
	.datab(!\E_iw[11]~q ),
	.datac(!\E_iw[16]~q ),
	.datad(!\E_iw[15]~q ),
	.datae(!\E_iw[13]~q ),
	.dataf(!\Equal209~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_rdctl~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_op_rdctl~0 .extended_lut = "off";
defparam \E_op_rdctl~0 .lut_mask = 64'hFFDFFFFFFFFFFFFF;
defparam \E_op_rdctl~0 .shared_arith = "off";

cyclonev_lcell_comb E_op_rdctl(
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_op_rdctl~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_rdctl~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_op_rdctl.extended_lut = "off";
defparam E_op_rdctl.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam E_op_rdctl.shared_arith = "off";

dffeas M_ctrl_rdctl_inst(
	.clk(clk_clk),
	.d(\E_op_rdctl~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_rdctl_inst~q ),
	.prn(vcc));
defparam M_ctrl_rdctl_inst.is_wysiwyg = "true";
defparam M_ctrl_rdctl_inst.power_up = "low";

cyclonev_lcell_comb \M_ctrl_mem_nxt~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[1]~q ),
	.datac(!\E_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ctrl_mem_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ctrl_mem_nxt~0 .extended_lut = "off";
defparam \M_ctrl_mem_nxt~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_ctrl_mem_nxt~0 .shared_arith = "off";

dffeas M_ctrl_mem(
	.clk(clk_clk),
	.d(\M_ctrl_mem_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_mem~q ),
	.prn(vcc));
defparam M_ctrl_mem.is_wysiwyg = "true";
defparam M_ctrl_mem.power_up = "low";

dffeas \A_inst_result[31] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.asdata(\M_alu_result[31]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[31]~q ),
	.prn(vcc));
defparam \A_inst_result[31] .is_wysiwyg = "true";
defparam \A_inst_result[31] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot~0 (
	.dataa(!\Equal171~0_combout ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_ctrl_shift_rot~0 .shared_arith = "off";

dffeas E_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_shift_rot~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot.is_wysiwyg = "true";
defparam E_ctrl_shift_rot.power_up = "low";

dffeas M_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\E_ctrl_shift_rot~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_shift_rot~q ),
	.prn(vcc));
defparam M_ctrl_shift_rot.is_wysiwyg = "true";
defparam M_ctrl_shift_rot.power_up = "low";

dffeas A_ctrl_shift_rot(
	.clk(clk_clk),
	.d(\M_ctrl_shift_rot~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_shift_rot~q ),
	.prn(vcc));
defparam A_ctrl_shift_rot.is_wysiwyg = "true";
defparam A_ctrl_shift_rot.power_up = "low";

cyclonev_lcell_comb \E_ld_bus~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[1]~q ),
	.datad(!\E_iw[4]~q ),
	.datae(!\E_iw[2]~q ),
	.dataf(!\Add17~37_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ld_bus~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ld_bus~0 .extended_lut = "off";
defparam \E_ld_bus~0 .lut_mask = 64'hFF7FFFFFFFFFFFFF;
defparam \E_ld_bus~0 .shared_arith = "off";

dffeas M_ctrl_ld_bypass(
	.clk(clk_clk),
	.d(\E_ld_bus~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_bypass~q ),
	.prn(vcc));
defparam M_ctrl_ld_bypass.is_wysiwyg = "true";
defparam M_ctrl_ld_bypass.power_up = "low";

dffeas A_ctrl_ld_bypass(
	.clk(clk_clk),
	.d(\M_ctrl_ld_bypass~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_ld_bypass~q ),
	.prn(vcc));
defparam A_ctrl_ld_bypass.is_wysiwyg = "true";
defparam A_ctrl_ld_bypass.power_up = "low";

cyclonev_lcell_comb \A_slow_inst_sel_nxt~0 (
	.dataa(!\A_dc_want_fill~q ),
	.datab(!\A_ctrl_ld_bypass~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_sel_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_sel_nxt~0 .extended_lut = "off";
defparam \A_slow_inst_sel_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \A_slow_inst_sel_nxt~0 .shared_arith = "off";

dffeas A_slow_inst_sel(
	.clk(clk_clk),
	.d(\A_slow_inst_sel_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_slow_inst_sel~q ),
	.prn(vcc));
defparam A_slow_inst_sel.is_wysiwyg = "true";
defparam A_slow_inst_sel.power_up = "low";

cyclonev_lcell_comb \E_ctrl_ld8_ld16~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[1]~q ),
	.datac(!\E_iw[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_ld8_ld16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_ld8_ld16~0 .extended_lut = "off";
defparam \E_ctrl_ld8_ld16~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \E_ctrl_ld8_ld16~0 .shared_arith = "off";

dffeas M_ctrl_ld8_ld16(
	.clk(clk_clk),
	.d(\E_ctrl_ld8_ld16~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld8_ld16~q ),
	.prn(vcc));
defparam M_ctrl_ld8_ld16.is_wysiwyg = "true";
defparam M_ctrl_ld8_ld16.power_up = "low";

dffeas A_ld_align_byte2_byte3_fill(
	.clk(clk_clk),
	.d(\M_ctrl_ld8_ld16~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ld_align_byte2_byte3_fill~q ),
	.prn(vcc));
defparam A_ld_align_byte2_byte3_fill.is_wysiwyg = "true";
defparam A_ld_align_byte2_byte3_fill.power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[29]~32 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_slow_inst_sel~q ),
	.datac(!\A_ld_align_byte2_byte3_fill~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[29]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[29]~32 .extended_lut = "off";
defparam \A_wr_data_unfiltered[29]~32 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \A_wr_data_unfiltered[29]~32 .shared_arith = "off";

dffeas \A_mul_partial_prod[31] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~57_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[31]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[31] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[31] .power_up = "low";

dffeas \A_mul_partial_prod[30] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~53_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[30]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[30] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[30] .power_up = "low";

dffeas \A_mul_partial_prod[29] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~49_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[29]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[29] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[29] .power_up = "low";

dffeas \A_mul_partial_prod[28] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~61_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[28]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[28] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[28] .power_up = "low";

dffeas \A_mul_partial_prod[27] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~25_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[27]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[27] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[27] .power_up = "low";

dffeas \A_mul_partial_prod[26] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~33_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[26]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[26] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[26] .power_up = "low";

dffeas \A_mul_partial_prod[25] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~9_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[25]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[25] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[25] .power_up = "low";

dffeas \A_mul_partial_prod[24] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~17_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[24]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[24] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[24] .power_up = "low";

dffeas \A_mul_partial_prod[23] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~41_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[23]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[23] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[23] .power_up = "low";

dffeas \A_mul_partial_prod[22] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~45_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[22]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[22] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[22] .power_up = "low";

dffeas \A_mul_partial_prod[21] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~1_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[21]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[21] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[21] .power_up = "low";

dffeas \A_mul_partial_prod[20] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~5_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[20]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[20] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[20] .power_up = "low";

dffeas \A_mul_partial_prod[19] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~29_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[19]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[19] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[19] .power_up = "low";

dffeas \A_mul_partial_prod[18] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~37_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[18]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[18] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[18] .power_up = "low";

dffeas \A_mul_partial_prod[17] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~13_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[17]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[17] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[17] .power_up = "low";

dffeas \A_mul_partial_prod[16] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|Add0~21_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[16]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[16] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[16] .power_up = "low";

dffeas \A_mul_partial_prod[15] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[15]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[15] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[15] .power_up = "low";

dffeas \A_mul_partial_prod[14] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[14]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[14] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[14] .power_up = "low";

dffeas \A_mul_partial_prod[13] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[13]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[13] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[13] .power_up = "low";

dffeas \A_mul_partial_prod[12] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[12]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[12] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[12] .power_up = "low";

dffeas \A_mul_partial_prod[11] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[11]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[11] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[11] .power_up = "low";

dffeas \A_mul_partial_prod[10] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[10]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[10] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[10] .power_up = "low";

dffeas \A_mul_partial_prod[9] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[9]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[9] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[9] .power_up = "low";

dffeas \A_mul_partial_prod[8] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[8]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[8] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[8] .power_up = "low";

dffeas \A_mul_partial_prod[7] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[7]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[7] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[7] .power_up = "low";

dffeas \A_mul_partial_prod[6] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[6]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[6] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[6] .power_up = "low";

dffeas \A_mul_partial_prod[5] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[5]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[5] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[5] .power_up = "low";

dffeas \A_mul_partial_prod[4] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[4]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[4] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[4] .power_up = "low";

dffeas \A_mul_partial_prod[3] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[3]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[3] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[3] .power_up = "low";

dffeas \A_mul_partial_prod[2] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[2]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[2] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[2] .power_up = "low";

dffeas \A_mul_partial_prod[1] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[1]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[1] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[1] .power_up = "low";

dffeas \A_mul_partial_prod[0] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_mult_cell|the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_partial_prod[0]~q ),
	.prn(vcc));
defparam \A_mul_partial_prod[0] .is_wysiwyg = "true";
defparam \A_mul_partial_prod[0] .power_up = "low";

cyclonev_lcell_comb \Add19~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[0]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~53_sumout ),
	.cout(\Add19~54 ),
	.shareout());
defparam \Add19~53 .extended_lut = "off";
defparam \Add19~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~53 .shared_arith = "off";

cyclonev_lcell_comb \always120~0 (
	.dataa(!\A_stall~combout ),
	.datab(!\M_valid_from_E~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always120~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always120~0 .extended_lut = "off";
defparam \always120~0 .lut_mask = 64'h7777777777777777;
defparam \always120~0 .shared_arith = "off";

cyclonev_lcell_comb \A_mul_cnt_nxt[0]~2 (
	.dataa(!\A_mul_stall~q ),
	.datab(!\A_mul_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mul_cnt_nxt[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mul_cnt_nxt[0]~2 .extended_lut = "off";
defparam \A_mul_cnt_nxt[0]~2 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \A_mul_cnt_nxt[0]~2 .shared_arith = "off";

dffeas \A_mul_cnt[0] (
	.clk(clk_clk),
	.d(\A_mul_cnt_nxt[0]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_cnt[0]~q ),
	.prn(vcc));
defparam \A_mul_cnt[0] .is_wysiwyg = "true";
defparam \A_mul_cnt[0] .power_up = "low";

cyclonev_lcell_comb \A_mul_cnt_nxt[1]~1 (
	.dataa(!\A_mul_stall~q ),
	.datab(!\A_mul_cnt[1]~q ),
	.datac(!\A_mul_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mul_cnt_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mul_cnt_nxt[1]~1 .extended_lut = "off";
defparam \A_mul_cnt_nxt[1]~1 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \A_mul_cnt_nxt[1]~1 .shared_arith = "off";

dffeas \A_mul_cnt[1] (
	.clk(clk_clk),
	.d(\A_mul_cnt_nxt[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_cnt[1]~q ),
	.prn(vcc));
defparam \A_mul_cnt[1] .is_wysiwyg = "true";
defparam \A_mul_cnt[1] .power_up = "low";

cyclonev_lcell_comb \A_mul_cnt_nxt[2]~0 (
	.dataa(!\A_mul_stall~q ),
	.datab(!\A_mul_cnt[2]~q ),
	.datac(!\A_mul_cnt[1]~q ),
	.datad(!\A_mul_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mul_cnt_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mul_cnt_nxt[2]~0 .extended_lut = "off";
defparam \A_mul_cnt_nxt[2]~0 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \A_mul_cnt_nxt[2]~0 .shared_arith = "off";

dffeas \A_mul_cnt[2] (
	.clk(clk_clk),
	.d(\A_mul_cnt_nxt[2]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_cnt[2]~q ),
	.prn(vcc));
defparam \A_mul_cnt[2] .is_wysiwyg = "true";
defparam \A_mul_cnt[2] .power_up = "low";

cyclonev_lcell_comb \A_mul_stall_nxt~0 (
	.dataa(!\A_mul_stall~q ),
	.datab(!\always120~0_combout ),
	.datac(!\M_ctrl_mul_lsw~q ),
	.datad(!\A_mul_cnt[2]~q ),
	.datae(!\A_mul_cnt[1]~q ),
	.dataf(!\A_mul_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mul_stall_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mul_stall_nxt~0 .extended_lut = "off";
defparam \A_mul_stall_nxt~0 .lut_mask = 64'hBFFFFFFF1FFFFFFF;
defparam \A_mul_stall_nxt~0 .shared_arith = "off";

dffeas A_mul_stall(
	.clk(clk_clk),
	.d(\A_mul_stall_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_stall~q ),
	.prn(vcc));
defparam A_mul_stall.is_wysiwyg = "true";
defparam A_mul_stall.power_up = "low";

dffeas A_mul_stall_d1(
	.clk(clk_clk),
	.d(\A_mul_stall~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_stall_d1~q ),
	.prn(vcc));
defparam A_mul_stall_d1.is_wysiwyg = "true";
defparam A_mul_stall_d1.power_up = "low";

dffeas A_mul_stall_d2(
	.clk(clk_clk),
	.d(\A_mul_stall_d1~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_stall_d2~q ),
	.prn(vcc));
defparam A_mul_stall_d2.is_wysiwyg = "true";
defparam A_mul_stall_d2.power_up = "low";

dffeas A_mul_stall_d3(
	.clk(clk_clk),
	.d(\A_mul_stall_d2~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mul_stall_d3~q ),
	.prn(vcc));
defparam A_mul_stall_d3.is_wysiwyg = "true";
defparam A_mul_stall_d3.power_up = "low";

dffeas \A_mul_result[0] (
	.clk(clk_clk),
	.d(\Add19~53_sumout ),
	.asdata(\A_mul_partial_prod[0]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[0]~q ),
	.prn(vcc));
defparam \A_mul_result[0] .is_wysiwyg = "true";
defparam \A_mul_result[0] .power_up = "low";

cyclonev_lcell_comb \Add19~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[1]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[1]~q ),
	.datag(gnd),
	.cin(\Add19~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~49_sumout ),
	.cout(\Add19~50 ),
	.shareout());
defparam \Add19~49 .extended_lut = "off";
defparam \Add19~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~49 .shared_arith = "off";

dffeas \A_mul_result[1] (
	.clk(clk_clk),
	.d(\Add19~49_sumout ),
	.asdata(\A_mul_partial_prod[1]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[1]~q ),
	.prn(vcc));
defparam \A_mul_result[1] .is_wysiwyg = "true";
defparam \A_mul_result[1] .power_up = "low";

cyclonev_lcell_comb \Add19~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[2]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[2]~q ),
	.datag(gnd),
	.cin(\Add19~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~1_sumout ),
	.cout(\Add19~2 ),
	.shareout());
defparam \Add19~1 .extended_lut = "off";
defparam \Add19~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~1 .shared_arith = "off";

dffeas \A_mul_result[2] (
	.clk(clk_clk),
	.d(\Add19~1_sumout ),
	.asdata(\A_mul_partial_prod[2]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[2]~q ),
	.prn(vcc));
defparam \A_mul_result[2] .is_wysiwyg = "true";
defparam \A_mul_result[2] .power_up = "low";

cyclonev_lcell_comb \Add19~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[3]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[3]~q ),
	.datag(gnd),
	.cin(\Add19~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~45_sumout ),
	.cout(\Add19~46 ),
	.shareout());
defparam \Add19~45 .extended_lut = "off";
defparam \Add19~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~45 .shared_arith = "off";

dffeas \A_mul_result[3] (
	.clk(clk_clk),
	.d(\Add19~45_sumout ),
	.asdata(\A_mul_partial_prod[3]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[3]~q ),
	.prn(vcc));
defparam \A_mul_result[3] .is_wysiwyg = "true";
defparam \A_mul_result[3] .power_up = "low";

cyclonev_lcell_comb \Add19~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[4]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[4]~q ),
	.datag(gnd),
	.cin(\Add19~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~41_sumout ),
	.cout(\Add19~42 ),
	.shareout());
defparam \Add19~41 .extended_lut = "off";
defparam \Add19~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~41 .shared_arith = "off";

dffeas \A_mul_result[4] (
	.clk(clk_clk),
	.d(\Add19~41_sumout ),
	.asdata(\A_mul_partial_prod[4]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[4]~q ),
	.prn(vcc));
defparam \A_mul_result[4] .is_wysiwyg = "true";
defparam \A_mul_result[4] .power_up = "low";

cyclonev_lcell_comb \Add19~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[5]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[5]~q ),
	.datag(gnd),
	.cin(\Add19~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~37_sumout ),
	.cout(\Add19~38 ),
	.shareout());
defparam \Add19~37 .extended_lut = "off";
defparam \Add19~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~37 .shared_arith = "off";

dffeas \A_mul_result[5] (
	.clk(clk_clk),
	.d(\Add19~37_sumout ),
	.asdata(\A_mul_partial_prod[5]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[5]~q ),
	.prn(vcc));
defparam \A_mul_result[5] .is_wysiwyg = "true";
defparam \A_mul_result[5] .power_up = "low";

cyclonev_lcell_comb \Add19~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[6]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[6]~q ),
	.datag(gnd),
	.cin(\Add19~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~33_sumout ),
	.cout(\Add19~34 ),
	.shareout());
defparam \Add19~33 .extended_lut = "off";
defparam \Add19~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~33 .shared_arith = "off";

dffeas \A_mul_result[6] (
	.clk(clk_clk),
	.d(\Add19~33_sumout ),
	.asdata(\A_mul_partial_prod[6]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[6]~q ),
	.prn(vcc));
defparam \A_mul_result[6] .is_wysiwyg = "true";
defparam \A_mul_result[6] .power_up = "low";

cyclonev_lcell_comb \Add19~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[7]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[7]~q ),
	.datag(gnd),
	.cin(\Add19~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~29_sumout ),
	.cout(\Add19~30 ),
	.shareout());
defparam \Add19~29 .extended_lut = "off";
defparam \Add19~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~29 .shared_arith = "off";

dffeas \A_mul_result[7] (
	.clk(clk_clk),
	.d(\Add19~29_sumout ),
	.asdata(\A_mul_partial_prod[7]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[7]~q ),
	.prn(vcc));
defparam \A_mul_result[7] .is_wysiwyg = "true";
defparam \A_mul_result[7] .power_up = "low";

cyclonev_lcell_comb \Add19~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[8]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[8]~q ),
	.datag(gnd),
	.cin(\Add19~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~25_sumout ),
	.cout(\Add19~26 ),
	.shareout());
defparam \Add19~25 .extended_lut = "off";
defparam \Add19~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~25 .shared_arith = "off";

dffeas \A_mul_result[8] (
	.clk(clk_clk),
	.d(\Add19~25_sumout ),
	.asdata(\A_mul_partial_prod[8]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[8]~q ),
	.prn(vcc));
defparam \A_mul_result[8] .is_wysiwyg = "true";
defparam \A_mul_result[8] .power_up = "low";

cyclonev_lcell_comb \Add19~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[9]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[9]~q ),
	.datag(gnd),
	.cin(\Add19~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~21_sumout ),
	.cout(\Add19~22 ),
	.shareout());
defparam \Add19~21 .extended_lut = "off";
defparam \Add19~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~21 .shared_arith = "off";

dffeas \A_mul_result[9] (
	.clk(clk_clk),
	.d(\Add19~21_sumout ),
	.asdata(\A_mul_partial_prod[9]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[9]~q ),
	.prn(vcc));
defparam \A_mul_result[9] .is_wysiwyg = "true";
defparam \A_mul_result[9] .power_up = "low";

cyclonev_lcell_comb \Add19~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[10]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[10]~q ),
	.datag(gnd),
	.cin(\Add19~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~17_sumout ),
	.cout(\Add19~18 ),
	.shareout());
defparam \Add19~17 .extended_lut = "off";
defparam \Add19~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~17 .shared_arith = "off";

dffeas \A_mul_result[10] (
	.clk(clk_clk),
	.d(\Add19~17_sumout ),
	.asdata(\A_mul_partial_prod[10]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[10]~q ),
	.prn(vcc));
defparam \A_mul_result[10] .is_wysiwyg = "true";
defparam \A_mul_result[10] .power_up = "low";

cyclonev_lcell_comb \Add19~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[11]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[11]~q ),
	.datag(gnd),
	.cin(\Add19~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~13_sumout ),
	.cout(\Add19~14 ),
	.shareout());
defparam \Add19~13 .extended_lut = "off";
defparam \Add19~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~13 .shared_arith = "off";

dffeas \A_mul_result[11] (
	.clk(clk_clk),
	.d(\Add19~13_sumout ),
	.asdata(\A_mul_partial_prod[11]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[11]~q ),
	.prn(vcc));
defparam \A_mul_result[11] .is_wysiwyg = "true";
defparam \A_mul_result[11] .power_up = "low";

cyclonev_lcell_comb \Add19~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[12]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[12]~q ),
	.datag(gnd),
	.cin(\Add19~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~9_sumout ),
	.cout(\Add19~10 ),
	.shareout());
defparam \Add19~9 .extended_lut = "off";
defparam \Add19~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~9 .shared_arith = "off";

dffeas \A_mul_result[12] (
	.clk(clk_clk),
	.d(\Add19~9_sumout ),
	.asdata(\A_mul_partial_prod[12]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[12]~q ),
	.prn(vcc));
defparam \A_mul_result[12] .is_wysiwyg = "true";
defparam \A_mul_result[12] .power_up = "low";

cyclonev_lcell_comb \Add19~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[13]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[13]~q ),
	.datag(gnd),
	.cin(\Add19~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~5_sumout ),
	.cout(\Add19~6 ),
	.shareout());
defparam \Add19~5 .extended_lut = "off";
defparam \Add19~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~5 .shared_arith = "off";

dffeas \A_mul_result[13] (
	.clk(clk_clk),
	.d(\Add19~5_sumout ),
	.asdata(\A_mul_partial_prod[13]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[13]~q ),
	.prn(vcc));
defparam \A_mul_result[13] .is_wysiwyg = "true";
defparam \A_mul_result[13] .power_up = "low";

cyclonev_lcell_comb \Add19~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[14]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[14]~q ),
	.datag(gnd),
	.cin(\Add19~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~109_sumout ),
	.cout(\Add19~110 ),
	.shareout());
defparam \Add19~109 .extended_lut = "off";
defparam \Add19~109 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~109 .shared_arith = "off";

dffeas \A_mul_result[14] (
	.clk(clk_clk),
	.d(\Add19~109_sumout ),
	.asdata(\A_mul_partial_prod[14]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[14]~q ),
	.prn(vcc));
defparam \A_mul_result[14] .is_wysiwyg = "true";
defparam \A_mul_result[14] .power_up = "low";

cyclonev_lcell_comb \Add19~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[15]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[15]~q ),
	.datag(gnd),
	.cin(\Add19~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~101_sumout ),
	.cout(\Add19~102 ),
	.shareout());
defparam \Add19~101 .extended_lut = "off";
defparam \Add19~101 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~101 .shared_arith = "off";

dffeas \A_mul_result[15] (
	.clk(clk_clk),
	.d(\Add19~101_sumout ),
	.asdata(\A_mul_partial_prod[15]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[15]~q ),
	.prn(vcc));
defparam \A_mul_result[15] .is_wysiwyg = "true";
defparam \A_mul_result[15] .power_up = "low";

cyclonev_lcell_comb \Add19~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[16]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[16]~q ),
	.datag(gnd),
	.cin(\Add19~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~77_sumout ),
	.cout(\Add19~78 ),
	.shareout());
defparam \Add19~77 .extended_lut = "off";
defparam \Add19~77 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~77 .shared_arith = "off";

dffeas \A_mul_result[16] (
	.clk(clk_clk),
	.d(\Add19~77_sumout ),
	.asdata(\A_mul_partial_prod[16]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[16]~q ),
	.prn(vcc));
defparam \A_mul_result[16] .is_wysiwyg = "true";
defparam \A_mul_result[16] .power_up = "low";

cyclonev_lcell_comb \Add19~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[17]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[17]~q ),
	.datag(gnd),
	.cin(\Add19~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~69_sumout ),
	.cout(\Add19~70 ),
	.shareout());
defparam \Add19~69 .extended_lut = "off";
defparam \Add19~69 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~69 .shared_arith = "off";

dffeas \A_mul_result[17] (
	.clk(clk_clk),
	.d(\Add19~69_sumout ),
	.asdata(\A_mul_partial_prod[17]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[17]~q ),
	.prn(vcc));
defparam \A_mul_result[17] .is_wysiwyg = "true";
defparam \A_mul_result[17] .power_up = "low";

cyclonev_lcell_comb \Add19~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[18]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[18]~q ),
	.datag(gnd),
	.cin(\Add19~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~93_sumout ),
	.cout(\Add19~94 ),
	.shareout());
defparam \Add19~93 .extended_lut = "off";
defparam \Add19~93 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~93 .shared_arith = "off";

dffeas \A_mul_result[18] (
	.clk(clk_clk),
	.d(\Add19~93_sumout ),
	.asdata(\A_mul_partial_prod[18]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[18]~q ),
	.prn(vcc));
defparam \A_mul_result[18] .is_wysiwyg = "true";
defparam \A_mul_result[18] .power_up = "low";

cyclonev_lcell_comb \Add19~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[19]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[19]~q ),
	.datag(gnd),
	.cin(\Add19~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~85_sumout ),
	.cout(\Add19~86 ),
	.shareout());
defparam \Add19~85 .extended_lut = "off";
defparam \Add19~85 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~85 .shared_arith = "off";

dffeas \A_mul_result[19] (
	.clk(clk_clk),
	.d(\Add19~85_sumout ),
	.asdata(\A_mul_partial_prod[19]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[19]~q ),
	.prn(vcc));
defparam \A_mul_result[19] .is_wysiwyg = "true";
defparam \A_mul_result[19] .power_up = "low";

cyclonev_lcell_comb \Add19~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[20]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[20]~q ),
	.datag(gnd),
	.cin(\Add19~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~61_sumout ),
	.cout(\Add19~62 ),
	.shareout());
defparam \Add19~61 .extended_lut = "off";
defparam \Add19~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~61 .shared_arith = "off";

dffeas \A_mul_result[20] (
	.clk(clk_clk),
	.d(\Add19~61_sumout ),
	.asdata(\A_mul_partial_prod[20]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[20]~q ),
	.prn(vcc));
defparam \A_mul_result[20] .is_wysiwyg = "true";
defparam \A_mul_result[20] .power_up = "low";

cyclonev_lcell_comb \Add19~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[21]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[21]~q ),
	.datag(gnd),
	.cin(\Add19~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~57_sumout ),
	.cout(\Add19~58 ),
	.shareout());
defparam \Add19~57 .extended_lut = "off";
defparam \Add19~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~57 .shared_arith = "off";

dffeas \A_mul_result[21] (
	.clk(clk_clk),
	.d(\Add19~57_sumout ),
	.asdata(\A_mul_partial_prod[21]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[21]~q ),
	.prn(vcc));
defparam \A_mul_result[21] .is_wysiwyg = "true";
defparam \A_mul_result[21] .power_up = "low";

cyclonev_lcell_comb \Add19~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[22]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[22]~q ),
	.datag(gnd),
	.cin(\Add19~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~105_sumout ),
	.cout(\Add19~106 ),
	.shareout());
defparam \Add19~105 .extended_lut = "off";
defparam \Add19~105 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~105 .shared_arith = "off";

dffeas \A_mul_result[22] (
	.clk(clk_clk),
	.d(\Add19~105_sumout ),
	.asdata(\A_mul_partial_prod[22]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[22]~q ),
	.prn(vcc));
defparam \A_mul_result[22] .is_wysiwyg = "true";
defparam \A_mul_result[22] .power_up = "low";

cyclonev_lcell_comb \Add19~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[23]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[23]~q ),
	.datag(gnd),
	.cin(\Add19~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~97_sumout ),
	.cout(\Add19~98 ),
	.shareout());
defparam \Add19~97 .extended_lut = "off";
defparam \Add19~97 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~97 .shared_arith = "off";

dffeas \A_mul_result[23] (
	.clk(clk_clk),
	.d(\Add19~97_sumout ),
	.asdata(\A_mul_partial_prod[23]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[23]~q ),
	.prn(vcc));
defparam \A_mul_result[23] .is_wysiwyg = "true";
defparam \A_mul_result[23] .power_up = "low";

cyclonev_lcell_comb \Add19~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[24]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[24]~q ),
	.datag(gnd),
	.cin(\Add19~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~73_sumout ),
	.cout(\Add19~74 ),
	.shareout());
defparam \Add19~73 .extended_lut = "off";
defparam \Add19~73 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~73 .shared_arith = "off";

dffeas \A_mul_result[24] (
	.clk(clk_clk),
	.d(\Add19~73_sumout ),
	.asdata(\A_mul_partial_prod[24]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[24]~q ),
	.prn(vcc));
defparam \A_mul_result[24] .is_wysiwyg = "true";
defparam \A_mul_result[24] .power_up = "low";

cyclonev_lcell_comb \Add19~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[25]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[25]~q ),
	.datag(gnd),
	.cin(\Add19~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~65_sumout ),
	.cout(\Add19~66 ),
	.shareout());
defparam \Add19~65 .extended_lut = "off";
defparam \Add19~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~65 .shared_arith = "off";

dffeas \A_mul_result[25] (
	.clk(clk_clk),
	.d(\Add19~65_sumout ),
	.asdata(\A_mul_partial_prod[25]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[25]~q ),
	.prn(vcc));
defparam \A_mul_result[25] .is_wysiwyg = "true";
defparam \A_mul_result[25] .power_up = "low";

cyclonev_lcell_comb \Add19~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[26]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[26]~q ),
	.datag(gnd),
	.cin(\Add19~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~89_sumout ),
	.cout(\Add19~90 ),
	.shareout());
defparam \Add19~89 .extended_lut = "off";
defparam \Add19~89 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~89 .shared_arith = "off";

dffeas \A_mul_result[26] (
	.clk(clk_clk),
	.d(\Add19~89_sumout ),
	.asdata(\A_mul_partial_prod[26]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[26]~q ),
	.prn(vcc));
defparam \A_mul_result[26] .is_wysiwyg = "true";
defparam \A_mul_result[26] .power_up = "low";

cyclonev_lcell_comb \Add19~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[27]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[27]~q ),
	.datag(gnd),
	.cin(\Add19~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~81_sumout ),
	.cout(\Add19~82 ),
	.shareout());
defparam \Add19~81 .extended_lut = "off";
defparam \Add19~81 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~81 .shared_arith = "off";

dffeas \A_mul_result[27] (
	.clk(clk_clk),
	.d(\Add19~81_sumout ),
	.asdata(\A_mul_partial_prod[27]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[27]~q ),
	.prn(vcc));
defparam \A_mul_result[27] .is_wysiwyg = "true";
defparam \A_mul_result[27] .power_up = "low";

cyclonev_lcell_comb \Add19~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[28]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[28]~q ),
	.datag(gnd),
	.cin(\Add19~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~125_sumout ),
	.cout(\Add19~126 ),
	.shareout());
defparam \Add19~125 .extended_lut = "off";
defparam \Add19~125 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~125 .shared_arith = "off";

dffeas \A_mul_result[28] (
	.clk(clk_clk),
	.d(\Add19~125_sumout ),
	.asdata(\A_mul_partial_prod[28]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[28]~q ),
	.prn(vcc));
defparam \A_mul_result[28] .is_wysiwyg = "true";
defparam \A_mul_result[28] .power_up = "low";

cyclonev_lcell_comb \Add19~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[29]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[29]~q ),
	.datag(gnd),
	.cin(\Add19~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~113_sumout ),
	.cout(\Add19~114 ),
	.shareout());
defparam \Add19~113 .extended_lut = "off";
defparam \Add19~113 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~113 .shared_arith = "off";

dffeas \A_mul_result[29] (
	.clk(clk_clk),
	.d(\Add19~113_sumout ),
	.asdata(\A_mul_partial_prod[29]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[29]~q ),
	.prn(vcc));
defparam \A_mul_result[29] .is_wysiwyg = "true";
defparam \A_mul_result[29] .power_up = "low";

cyclonev_lcell_comb \Add19~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[30]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[30]~q ),
	.datag(gnd),
	.cin(\Add19~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~117_sumout ),
	.cout(\Add19~118 ),
	.shareout());
defparam \Add19~117 .extended_lut = "off";
defparam \Add19~117 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~117 .shared_arith = "off";

dffeas \A_mul_result[30] (
	.clk(clk_clk),
	.d(\Add19~117_sumout ),
	.asdata(\A_mul_partial_prod[30]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[30]~q ),
	.prn(vcc));
defparam \A_mul_result[30] .is_wysiwyg = "true";
defparam \A_mul_result[30] .power_up = "low";

cyclonev_lcell_comb \Add19~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\A_mul_result[31]~q ),
	.datae(gnd),
	.dataf(!\A_mul_partial_prod[31]~q ),
	.datag(gnd),
	.cin(\Add19~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add19~121_sumout ),
	.cout(),
	.shareout());
defparam \Add19~121 .extended_lut = "off";
defparam \Add19~121 .lut_mask = 64'h0000FF00000000FF;
defparam \Add19~121 .shared_arith = "off";

dffeas \A_mul_result[31] (
	.clk(clk_clk),
	.d(\Add19~121_sumout ),
	.asdata(\A_mul_partial_prod[31]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_mul_stall_d3~q ),
	.ena(vcc),
	.q(\A_mul_result[31]~q ),
	.prn(vcc));
defparam \A_mul_result[31] .is_wysiwyg = "true";
defparam \A_mul_result[31] .power_up = "low";

dffeas \D_iw[6] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[6]~q ),
	.prn(vcc));
defparam \D_iw[6] .is_wysiwyg = "true";
defparam \D_iw[6] .power_up = "low";

dffeas \E_compare_op[0] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[0]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_compare_op[0]~q ),
	.prn(vcc));
defparam \E_compare_op[0] .is_wysiwyg = "true";
defparam \E_compare_op[0] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[0]~28 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(gnd),
	.datad(!\Equal297~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~28 .extended_lut = "off";
defparam \D_src2_reg[0]~28 .lut_mask = 64'hFFBBFFBBFFBBFFBB;
defparam \D_src2_reg[0]~28 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~20 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[27]~6_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~20 .extended_lut = "off";
defparam \E_alu_result~20 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~20 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[27] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~20_combout ),
	.datac(!\Add17~97_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[27]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[27] .extended_lut = "off";
defparam \E_alu_result[27] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[27] .shared_arith = "off";

dffeas \M_alu_result[27] (
	.clk(clk_clk),
	.d(\E_alu_result[27]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[27]~q ),
	.prn(vcc));
defparam \M_alu_result[27] .is_wysiwyg = "true";
defparam \M_alu_result[27] .power_up = "low";

dffeas \A_inst_result[27] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[27] ),
	.asdata(\M_alu_result[27]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[27]~q ),
	.prn(vcc));
defparam \A_inst_result[27] .is_wysiwyg = "true";
defparam \A_inst_result[27] .power_up = "low";

cyclonev_lcell_comb \E_ctrl_ld_signed~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[1]~q ),
	.datac(!\E_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_ld_signed~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_ld_signed~0 .extended_lut = "off";
defparam \E_ctrl_ld_signed~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_ctrl_ld_signed~0 .shared_arith = "off";

dffeas M_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\E_ctrl_ld_signed~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_signed~q ),
	.prn(vcc));
defparam M_ctrl_ld_signed.is_wysiwyg = "true";
defparam M_ctrl_ld_signed.power_up = "low";

dffeas A_ctrl_ld_signed(
	.clk(clk_clk),
	.d(\M_ctrl_ld_signed~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_ld_signed~q ),
	.prn(vcc));
defparam A_ctrl_ld_signed.is_wysiwyg = "true";
defparam A_ctrl_ld_signed.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_right_arith~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\Equal171~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_right_arith~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_right_arith~0 .extended_lut = "off";
defparam \D_ctrl_shift_right_arith~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \D_ctrl_shift_right_arith~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_right_arith~1 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_ctrl_shift_right_arith~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_right_arith~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_right_arith~1 .extended_lut = "off";
defparam \D_ctrl_shift_right_arith~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \D_ctrl_shift_right_arith~1 .shared_arith = "off";

dffeas E_ctrl_shift_right_arith(
	.clk(clk_clk),
	.d(\D_ctrl_shift_right_arith~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_shift_right_arith~q ),
	.prn(vcc));
defparam E_ctrl_shift_right_arith.is_wysiwyg = "true";
defparam E_ctrl_shift_right_arith.power_up = "low";

cyclonev_lcell_comb \E_rot_fill_bit~0 (
	.dataa(!\E_src1[31]~q ),
	.datab(!\E_ctrl_shift_right_arith~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_fill_bit~0 .extended_lut = "off";
defparam \E_rot_fill_bit~0 .lut_mask = 64'h7777777777777777;
defparam \E_rot_fill_bit~0 .shared_arith = "off";

dffeas M_rot_fill_bit(
	.clk(clk_clk),
	.d(\E_rot_fill_bit~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_fill_bit~q ),
	.prn(vcc));
defparam M_rot_fill_bit.is_wysiwyg = "true";
defparam M_rot_fill_bit.power_up = "low";

dffeas \D_iw[8] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[8]~q ),
	.prn(vcc));
defparam \D_iw[8] .is_wysiwyg = "true";
defparam \D_iw[8] .power_up = "low";

dffeas \d_readdata_d1[2] (
	.clk(clk_clk),
	.d(d_readdata[2]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[2]~q ),
	.prn(vcc));
defparam \d_readdata_d1[2] .is_wysiwyg = "true";
defparam \d_readdata_d1[2] .power_up = "low";

dffeas \d_readdata_d1[10] (
	.clk(clk_clk),
	.d(d_readdata[10]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[10]~q ),
	.prn(vcc));
defparam \d_readdata_d1[10] .is_wysiwyg = "true";
defparam \d_readdata_d1[10] .power_up = "low";

dffeas \d_readdata_d1[18] (
	.clk(clk_clk),
	.d(d_readdata[18]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[18]~q ),
	.prn(vcc));
defparam \d_readdata_d1[18] .is_wysiwyg = "true";
defparam \d_readdata_d1[18] .power_up = "low";

dffeas \d_readdata_d1[26] (
	.clk(clk_clk),
	.d(d_readdata[26]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[26]~q ),
	.prn(vcc));
defparam \d_readdata_d1[26] .is_wysiwyg = "true";
defparam \d_readdata_d1[26] .power_up = "low";

dffeas \M_alu_result[0] (
	.clk(clk_clk),
	.d(\E_alu_result[0]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[0]~q ),
	.prn(vcc));
defparam \M_alu_result[0] .is_wysiwyg = "true";
defparam \M_alu_result[0] .power_up = "low";

cyclonev_lcell_comb \Equal184~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_ctrl_ld8_ld16~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal184~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal184~0 .extended_lut = "off";
defparam \Equal184~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal184~0 .shared_arith = "off";

dffeas M_ctrl_ld8(
	.clk(clk_clk),
	.d(\Equal184~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld8~q ),
	.prn(vcc));
defparam M_ctrl_ld8.is_wysiwyg = "true";
defparam M_ctrl_ld8.power_up = "low";

cyclonev_lcell_comb \M_ld_align_sh8~0 (
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\M_ctrl_ld8~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ld_align_sh8~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ld_align_sh8~0 .extended_lut = "off";
defparam \M_ld_align_sh8~0 .lut_mask = 64'h7777777777777777;
defparam \M_ld_align_sh8~0 .shared_arith = "off";

dffeas A_ld_align_sh8(
	.clk(clk_clk),
	.d(\M_ld_align_sh8~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ld_align_sh8~q ),
	.prn(vcc));
defparam A_ld_align_sh8.is_wysiwyg = "true";
defparam A_ld_align_sh8.power_up = "low";

dffeas \D_iw[7] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[7]~q ),
	.prn(vcc));
defparam \D_iw[7] .is_wysiwyg = "true";
defparam \D_iw[7] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[5]~3 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\M_regnum_b_cmp_D~q ),
	.datac(!\A_regnum_b_cmp_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~3 .extended_lut = "off";
defparam \D_src2_reg[5]~3 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \D_src2_reg[5]~3 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[5]~4 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\M_regnum_b_cmp_D~q ),
	.datac(!\A_regnum_b_cmp_D~q ),
	.datad(!\W_regnum_b_cmp_D~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~4 .extended_lut = "off";
defparam \D_src2_reg[5]~4 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \D_src2_reg[5]~4 .shared_arith = "off";

dffeas \d_readdata_d1[1] (
	.clk(clk_clk),
	.d(d_readdata[1]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[1]~q ),
	.prn(vcc));
defparam \d_readdata_d1[1] .is_wysiwyg = "true";
defparam \d_readdata_d1[1] .power_up = "low";

dffeas \d_readdata_d1[9] (
	.clk(clk_clk),
	.d(d_readdata[9]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[9]~q ),
	.prn(vcc));
defparam \d_readdata_d1[9] .is_wysiwyg = "true";
defparam \d_readdata_d1[9] .power_up = "low";

dffeas \d_readdata_d1[17] (
	.clk(clk_clk),
	.d(d_readdata[17]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[17]~q ),
	.prn(vcc));
defparam \d_readdata_d1[17] .is_wysiwyg = "true";
defparam \d_readdata_d1[17] .power_up = "low";

dffeas \d_readdata_d1[25] (
	.clk(clk_clk),
	.d(d_readdata[25]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[25]~q ),
	.prn(vcc));
defparam \d_readdata_d1[25] .is_wysiwyg = "true";
defparam \d_readdata_d1[25] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte0_data_aligned_nxt[1]~6 (
	.dataa(!\d_readdata_d1[1]~q ),
	.datab(!\d_readdata_d1[9]~q ),
	.datac(!\d_readdata_d1[17]~q ),
	.datad(!\d_readdata_d1[25]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte0_data_aligned_nxt[1]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte0_data_aligned_nxt[1]~6 .extended_lut = "off";
defparam \A_slow_ld_byte0_data_aligned_nxt[1]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_ld_byte0_data_aligned_nxt[1]~6 .shared_arith = "off";

dffeas d_readdatavalid_d1(
	.clk(clk_clk),
	.d(d_readdatavalid),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdatavalid_d1~q ),
	.prn(vcc));
defparam d_readdatavalid_d1.is_wysiwyg = "true";
defparam d_readdatavalid_d1.power_up = "low";

dffeas \D_iw[10] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[10]~q ),
	.prn(vcc));
defparam \D_iw[10] .is_wysiwyg = "true";
defparam \D_iw[10] .power_up = "low";

dffeas \d_readdata_d1[4] (
	.clk(clk_clk),
	.d(d_readdata[4]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[4]~q ),
	.prn(vcc));
defparam \d_readdata_d1[4] .is_wysiwyg = "true";
defparam \d_readdata_d1[4] .power_up = "low";

dffeas \d_readdata_d1[12] (
	.clk(clk_clk),
	.d(d_readdata[12]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[12]~q ),
	.prn(vcc));
defparam \d_readdata_d1[12] .is_wysiwyg = "true";
defparam \d_readdata_d1[12] .power_up = "low";

dffeas \d_readdata_d1[20] (
	.clk(clk_clk),
	.d(d_readdata[20]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[20]~q ),
	.prn(vcc));
defparam \d_readdata_d1[20] .is_wysiwyg = "true";
defparam \d_readdata_d1[20] .power_up = "low";

dffeas \d_readdata_d1[28] (
	.clk(clk_clk),
	.d(d_readdata[28]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[28]~q ),
	.prn(vcc));
defparam \d_readdata_d1[28] .is_wysiwyg = "true";
defparam \d_readdata_d1[28] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte0_data_aligned_nxt[4]~4 (
	.dataa(!\d_readdata_d1[4]~q ),
	.datab(!\d_readdata_d1[12]~q ),
	.datac(!\d_readdata_d1[20]~q ),
	.datad(!\d_readdata_d1[28]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte0_data_aligned_nxt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte0_data_aligned_nxt[4]~4 .extended_lut = "off";
defparam \A_slow_ld_byte0_data_aligned_nxt[4]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_ld_byte0_data_aligned_nxt[4]~4 .shared_arith = "off";

dffeas \A_slow_inst_result[4] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte0_data_aligned_nxt[4]~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[4]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[4] .is_wysiwyg = "true";
defparam \A_slow_inst_result[4] .power_up = "low";

dffeas \A_inst_result[4] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[4] ),
	.asdata(\M_alu_result[4]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[4]~q ),
	.prn(vcc));
defparam \A_inst_result[4] .is_wysiwyg = "true";
defparam \A_inst_result[4] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[13]~8 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[13]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[13]~8 .extended_lut = "off";
defparam \D_src2_reg[13]~8 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \D_src2_reg[13]~8 .shared_arith = "off";

dffeas \D_iw[9] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[9]~q ),
	.prn(vcc));
defparam \D_iw[9] .is_wysiwyg = "true";
defparam \D_iw[9] .power_up = "low";

dffeas \d_readdata_d1[3] (
	.clk(clk_clk),
	.d(d_readdata[3]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[3]~q ),
	.prn(vcc));
defparam \d_readdata_d1[3] .is_wysiwyg = "true";
defparam \d_readdata_d1[3] .power_up = "low";

dffeas \d_readdata_d1[11] (
	.clk(clk_clk),
	.d(d_readdata[11]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[11]~q ),
	.prn(vcc));
defparam \d_readdata_d1[11] .is_wysiwyg = "true";
defparam \d_readdata_d1[11] .power_up = "low";

dffeas \d_readdata_d1[19] (
	.clk(clk_clk),
	.d(d_readdata[19]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[19]~q ),
	.prn(vcc));
defparam \d_readdata_d1[19] .is_wysiwyg = "true";
defparam \d_readdata_d1[19] .power_up = "low";

dffeas \d_readdata_d1[27] (
	.clk(clk_clk),
	.d(d_readdata[27]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[27]~q ),
	.prn(vcc));
defparam \d_readdata_d1[27] .is_wysiwyg = "true";
defparam \d_readdata_d1[27] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte0_data_aligned_nxt[3]~5 (
	.dataa(!\d_readdata_d1[3]~q ),
	.datab(!\d_readdata_d1[11]~q ),
	.datac(!\d_readdata_d1[19]~q ),
	.datad(!\d_readdata_d1[27]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte0_data_aligned_nxt[3]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte0_data_aligned_nxt[3]~5 .extended_lut = "off";
defparam \A_slow_ld_byte0_data_aligned_nxt[3]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_ld_byte0_data_aligned_nxt[3]~5 .shared_arith = "off";

dffeas \A_slow_inst_result[3] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte0_data_aligned_nxt[3]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[3]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[3] .is_wysiwyg = "true";
defparam \A_slow_inst_result[3] .power_up = "low";

dffeas \A_inst_result[3] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[3] ),
	.asdata(\M_alu_result[3]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[3]~q ),
	.prn(vcc));
defparam \A_inst_result[3] .is_wysiwyg = "true";
defparam \A_inst_result[3] .power_up = "low";

dffeas E_ctrl_shift_rot_right(
	.clk(clk_clk),
	.d(\D_ctrl_shift_right_arith~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_shift_rot_right~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot_right.is_wysiwyg = "true";
defparam E_ctrl_shift_rot_right.power_up = "low";

cyclonev_lcell_comb \D_ctrl_shift_rot_left~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\Equal171~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot_left~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot_left~0 .extended_lut = "off";
defparam \D_ctrl_shift_rot_left~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \D_ctrl_shift_rot_left~0 .shared_arith = "off";

dffeas E_ctrl_shift_rot_left(
	.clk(clk_clk),
	.d(\D_ctrl_shift_rot_left~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_shift_rot_left~q ),
	.prn(vcc));
defparam E_ctrl_shift_rot_left.is_wysiwyg = "true";
defparam E_ctrl_shift_rot_left.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill1~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(!\E_ctrl_shift_rot_left~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill1~0 .extended_lut = "off";
defparam \E_rot_sel_fill1~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_sel_fill1~0 .shared_arith = "off";

dffeas M_rot_sel_fill1(
	.clk(clk_clk),
	.d(\E_rot_sel_fill1~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_sel_fill1~q ),
	.prn(vcc));
defparam M_rot_sel_fill1.is_wysiwyg = "true";
defparam M_rot_sel_fill1.power_up = "low";

dffeas \d_readdata_d1[7] (
	.clk(clk_clk),
	.d(d_readdata[7]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[7]~q ),
	.prn(vcc));
defparam \d_readdata_d1[7] .is_wysiwyg = "true";
defparam \d_readdata_d1[7] .power_up = "low";

dffeas \d_readdata_d1[15] (
	.clk(clk_clk),
	.d(d_readdata[15]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[15]~q ),
	.prn(vcc));
defparam \d_readdata_d1[15] .is_wysiwyg = "true";
defparam \d_readdata_d1[15] .power_up = "low";

dffeas \d_readdata_d1[23] (
	.clk(clk_clk),
	.d(d_readdata[23]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[23]~q ),
	.prn(vcc));
defparam \d_readdata_d1[23] .is_wysiwyg = "true";
defparam \d_readdata_d1[23] .power_up = "low";

dffeas \d_readdata_d1[31] (
	.clk(clk_clk),
	.d(d_readdata[31]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[31]~q ),
	.prn(vcc));
defparam \d_readdata_d1[31] .is_wysiwyg = "true";
defparam \d_readdata_d1[31] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte0_data_aligned_nxt[7]~1 (
	.dataa(!\d_readdata_d1[7]~q ),
	.datab(!\d_readdata_d1[15]~q ),
	.datac(!\d_readdata_d1[23]~q ),
	.datad(!\d_readdata_d1[31]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte0_data_aligned_nxt[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte0_data_aligned_nxt[7]~1 .extended_lut = "off";
defparam \A_slow_ld_byte0_data_aligned_nxt[7]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_ld_byte0_data_aligned_nxt[7]~1 .shared_arith = "off";

dffeas \A_slow_inst_result[7] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte0_data_aligned_nxt[7]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[7]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[7] .is_wysiwyg = "true";
defparam \A_slow_inst_result[7] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[7]~14 (
	.dataa(!\M_alu_result[7]~q ),
	.datab(!\D_src2_reg[5]~3_combout ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\W_wr_data[7]~q ),
	.datae(!\A_wr_data_unfiltered[7]~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[7]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[7]~14 .extended_lut = "off";
defparam \D_src2_reg[7]~14 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[7]~14 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[7]~15 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_src2_reg[7]~14_combout ),
	.datad(!\E_alu_result[7]~combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[7] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[7]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[7]~15 .extended_lut = "off";
defparam \D_src2_reg[7]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[7]~15 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_hi_imm16~0 (
	.dataa(!\F_iw[5]~1_combout ),
	.datab(!\F_iw[2]~5_combout ),
	.datac(!\F_iw[0]~9_combout ),
	.datad(!\F_iw[1]~3_combout ),
	.datae(!\F_iw[4]~4_combout ),
	.dataf(!\F_iw[3]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_hi_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_hi_imm16~0 .extended_lut = "off";
defparam \F_ctrl_hi_imm16~0 .lut_mask = 64'hFFF7FFFFFFFFFFFF;
defparam \F_ctrl_hi_imm16~0 .shared_arith = "off";

dffeas D_ctrl_hi_imm16(
	.clk(clk_clk),
	.d(\F_ctrl_hi_imm16~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_hi_imm16~q ),
	.prn(vcc));
defparam D_ctrl_hi_imm16.is_wysiwyg = "true";
defparam D_ctrl_hi_imm16.power_up = "low";

cyclonev_lcell_comb \E_src2[14]~0 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_ctrl_src2_choose_imm~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src2[14]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src2[14]~0 .extended_lut = "off";
defparam \E_src2[14]~0 .lut_mask = 64'h7777777777777777;
defparam \E_src2[14]~0 .shared_arith = "off";

dffeas \E_src2[7] (
	.clk(clk_clk),
	.d(\D_iw[13]~q ),
	.asdata(\D_src2_reg[7]~15_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[7]~q ),
	.prn(vcc));
defparam \E_src2[7] .is_wysiwyg = "true";
defparam \E_src2[7] .power_up = "low";

dffeas \d_readdata_d1[6] (
	.clk(clk_clk),
	.d(d_readdata[6]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[6]~q ),
	.prn(vcc));
defparam \d_readdata_d1[6] .is_wysiwyg = "true";
defparam \d_readdata_d1[6] .power_up = "low";

dffeas \d_readdata_d1[14] (
	.clk(clk_clk),
	.d(d_readdata[14]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[14]~q ),
	.prn(vcc));
defparam \d_readdata_d1[14] .is_wysiwyg = "true";
defparam \d_readdata_d1[14] .power_up = "low";

dffeas \d_readdata_d1[22] (
	.clk(clk_clk),
	.d(d_readdata[22]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[22]~q ),
	.prn(vcc));
defparam \d_readdata_d1[22] .is_wysiwyg = "true";
defparam \d_readdata_d1[22] .power_up = "low";

dffeas \d_readdata_d1[30] (
	.clk(clk_clk),
	.d(d_readdata[30]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[30]~q ),
	.prn(vcc));
defparam \d_readdata_d1[30] .is_wysiwyg = "true";
defparam \d_readdata_d1[30] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte0_data_aligned_nxt[6]~2 (
	.dataa(!\d_readdata_d1[6]~q ),
	.datab(!\d_readdata_d1[14]~q ),
	.datac(!\d_readdata_d1[22]~q ),
	.datad(!\d_readdata_d1[30]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte0_data_aligned_nxt[6]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte0_data_aligned_nxt[6]~2 .extended_lut = "off";
defparam \A_slow_ld_byte0_data_aligned_nxt[6]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_ld_byte0_data_aligned_nxt[6]~2 .shared_arith = "off";

dffeas \A_slow_inst_result[6] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte0_data_aligned_nxt[6]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[6]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[6] .is_wysiwyg = "true";
defparam \A_slow_inst_result[6] .power_up = "low";

dffeas \A_inst_result[6] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[6] ),
	.asdata(\M_alu_result[6]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[6]~q ),
	.prn(vcc));
defparam \A_inst_result[6] .is_wysiwyg = "true";
defparam \A_inst_result[6] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[6]~7 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[6]~7 .extended_lut = "off";
defparam \E_rot_mask[6]~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[6]~7 .shared_arith = "off";

dffeas \M_rot_mask[6] (
	.clk(clk_clk),
	.d(\E_rot_mask[6]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[6]~q ),
	.prn(vcc));
defparam \M_rot_mask[6] .is_wysiwyg = "true";
defparam \M_rot_mask[6] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[2]~0 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[2]~0 .extended_lut = "off";
defparam \E_rot_mask[2]~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[2]~0 .shared_arith = "off";

dffeas \M_rot_mask[2] (
	.clk(clk_clk),
	.d(\E_rot_mask[2]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[2]~q ),
	.prn(vcc));
defparam \M_rot_mask[2] .is_wysiwyg = "true";
defparam \M_rot_mask[2] .power_up = "low";

dffeas \d_readdata_d1[5] (
	.clk(clk_clk),
	.d(d_readdata[5]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[5]~q ),
	.prn(vcc));
defparam \d_readdata_d1[5] .is_wysiwyg = "true";
defparam \d_readdata_d1[5] .power_up = "low";

dffeas \d_readdata_d1[13] (
	.clk(clk_clk),
	.d(d_readdata[13]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[13]~q ),
	.prn(vcc));
defparam \d_readdata_d1[13] .is_wysiwyg = "true";
defparam \d_readdata_d1[13] .power_up = "low";

dffeas \d_readdata_d1[21] (
	.clk(clk_clk),
	.d(d_readdata[21]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[21]~q ),
	.prn(vcc));
defparam \d_readdata_d1[21] .is_wysiwyg = "true";
defparam \d_readdata_d1[21] .power_up = "low";

dffeas \d_readdata_d1[29] (
	.clk(clk_clk),
	.d(d_readdata[29]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[29]~q ),
	.prn(vcc));
defparam \d_readdata_d1[29] .is_wysiwyg = "true";
defparam \d_readdata_d1[29] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte0_data_aligned_nxt[5]~3 (
	.dataa(!\d_readdata_d1[5]~q ),
	.datab(!\d_readdata_d1[13]~q ),
	.datac(!\d_readdata_d1[21]~q ),
	.datad(!\d_readdata_d1[29]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte0_data_aligned_nxt[5]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte0_data_aligned_nxt[5]~3 .extended_lut = "off";
defparam \A_slow_ld_byte0_data_aligned_nxt[5]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_ld_byte0_data_aligned_nxt[5]~3 .shared_arith = "off";

dffeas \A_slow_inst_result[5] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte0_data_aligned_nxt[5]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[5]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[5] .is_wysiwyg = "true";
defparam \A_slow_inst_result[5] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[5]~18 (
	.dataa(!\M_alu_result[5]~q ),
	.datab(!\D_src2_reg[5]~3_combout ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\W_wr_data[5]~q ),
	.datae(!\A_wr_data_unfiltered[5]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~18 .extended_lut = "off";
defparam \D_src2_reg[5]~18 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[5]~18 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[5]~19 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_src2_reg[5]~18_combout ),
	.datad(!\E_alu_result[5]~combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[5] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[5]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[5]~19 .extended_lut = "off";
defparam \D_src2_reg[5]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[5]~19 .shared_arith = "off";

dffeas \E_src2[5] (
	.clk(clk_clk),
	.d(\D_iw[11]~q ),
	.asdata(\D_src2_reg[5]~19_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[5]~q ),
	.prn(vcc));
defparam \E_src2[5] .is_wysiwyg = "true";
defparam \E_src2[5] .power_up = "low";

cyclonev_lcell_comb \E_regnum_a_cmp_F~0 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datac(!\E_dst_regnum[0]~q ),
	.datad(!\E_dst_regnum[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \E_regnum_a_cmp_F~0 .lut_mask = 64'h6996699669966996;
defparam \E_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \E_regnum_a_cmp_F~1 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datac(!\E_dst_regnum[3]~q ),
	.datad(!\E_dst_regnum[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_a_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_a_cmp_F~1 .extended_lut = "off";
defparam \E_regnum_a_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \E_regnum_a_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb E_regnum_a_cmp_F(
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datab(!\E_dst_regnum[2]~q ),
	.datac(!\E_wr_dst_reg~0_combout ),
	.datad(!\E_regnum_a_cmp_F~0_combout ),
	.datae(!\E_regnum_a_cmp_F~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_regnum_a_cmp_F.extended_lut = "off";
defparam E_regnum_a_cmp_F.lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam E_regnum_a_cmp_F.shared_arith = "off";

cyclonev_lcell_comb \D_regnum_a_cmp_F~0 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datab(!\D_dst_regnum[0]~2_combout ),
	.datac(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datad(!\D_dst_regnum[2]~3_combout ),
	.datae(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(!\D_dst_regnum[3]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \D_regnum_a_cmp_F~0 .lut_mask = 64'h6996966996696996;
defparam \D_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb D_regnum_a_cmp_F(
	.dataa(!\D_dst_regnum[1]~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datac(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datad(!\D_dst_regnum[4]~1_combout ),
	.datae(!\D_wr_dst_reg~combout ),
	.dataf(!\D_regnum_a_cmp_F~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_regnum_a_cmp_F.extended_lut = "off";
defparam D_regnum_a_cmp_F.lut_mask = 64'h6996FFFFFFFFFFFF;
defparam D_regnum_a_cmp_F.shared_arith = "off";

dffeas E_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\D_regnum_a_cmp_F~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_stall~combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam E_regnum_a_cmp_D.is_wysiwyg = "true";
defparam E_regnum_a_cmp_D.power_up = "low";

dffeas M_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\E_regnum_a_cmp_F~combout ),
	.asdata(\E_regnum_a_cmp_D~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(\A_stall~combout ),
	.q(\M_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam M_regnum_a_cmp_D.is_wysiwyg = "true";
defparam M_regnum_a_cmp_D.power_up = "low";

cyclonev_lcell_comb \A_regnum_a_cmp_F~0 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datac(!\A_wr_dst_reg_from_M~q ),
	.datad(!\A_dst_regnum_from_M[0]~q ),
	.datae(!\A_dst_regnum_from_M[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \A_regnum_a_cmp_F~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \A_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \A_regnum_a_cmp_F~1 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datac(!\A_dst_regnum_from_M[2]~q ),
	.datad(!\A_dst_regnum_from_M[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_a_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_regnum_a_cmp_F~1 .extended_lut = "off";
defparam \A_regnum_a_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \A_regnum_a_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb A_regnum_a_cmp_F(
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datab(!\A_dst_regnum_from_M[4]~q ),
	.datac(!\A_regnum_a_cmp_F~0_combout ),
	.datad(!\A_regnum_a_cmp_F~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_regnum_a_cmp_F.extended_lut = "off";
defparam A_regnum_a_cmp_F.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam A_regnum_a_cmp_F.shared_arith = "off";

cyclonev_lcell_comb \M_regnum_a_cmp_F~0 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.datac(!\M_wr_dst_reg_from_E~q ),
	.datad(!\M_dst_regnum[0]~q ),
	.datae(!\M_dst_regnum[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_a_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_a_cmp_F~0 .extended_lut = "off";
defparam \M_regnum_a_cmp_F~0 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \M_regnum_a_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \M_regnum_a_cmp_F~1 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.datac(!\M_dst_regnum[2]~q ),
	.datad(!\M_dst_regnum[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_a_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_regnum_a_cmp_F~1 .extended_lut = "off";
defparam \M_regnum_a_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \M_regnum_a_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb M_regnum_a_cmp_F(
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.datab(!\M_dst_regnum[4]~q ),
	.datac(!\M_regnum_a_cmp_F~0_combout ),
	.datad(!\M_regnum_a_cmp_F~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_regnum_a_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_regnum_a_cmp_F.extended_lut = "off";
defparam M_regnum_a_cmp_F.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam M_regnum_a_cmp_F.shared_arith = "off";

dffeas A_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\M_regnum_a_cmp_F~combout ),
	.asdata(\M_regnum_a_cmp_D~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(\A_stall~combout ),
	.q(\A_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam A_regnum_a_cmp_D.is_wysiwyg = "true";
defparam A_regnum_a_cmp_D.power_up = "low";

dffeas W_regnum_a_cmp_D(
	.clk(clk_clk),
	.d(\A_regnum_a_cmp_F~combout ),
	.asdata(\A_regnum_a_cmp_D~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(vcc),
	.q(\W_regnum_a_cmp_D~q ),
	.prn(vcc));
defparam W_regnum_a_cmp_D.is_wysiwyg = "true";
defparam W_regnum_a_cmp_D.power_up = "low";

cyclonev_lcell_comb \E_src1[7]~0 (
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\M_regnum_a_cmp_D~q ),
	.datac(!\W_regnum_a_cmp_D~q ),
	.datad(!\A_regnum_a_cmp_D~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[7]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[7]~0 .extended_lut = "off";
defparam \E_src1[7]~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \E_src1[7]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_src1[7]~1 (
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\M_regnum_a_cmp_D~q ),
	.datac(!\A_regnum_a_cmp_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src1[7]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src1[7]~1 .extended_lut = "off";
defparam \E_src1[7]~1 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_src1[7]~1 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_reg[4]~10 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[4] ),
	.datab(!\W_wr_data[4]~q ),
	.datac(!\M_alu_result[4]~q ),
	.datad(!\A_wr_data_unfiltered[4]~25_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[4]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[4]~10 .extended_lut = "off";
defparam \D_src1_reg[4]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[4]~10 .shared_arith = "off";

dffeas \D_iw[28] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[28] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[28]~q ),
	.prn(vcc));
defparam \D_iw[28] .is_wysiwyg = "true";
defparam \D_iw[28] .power_up = "low";

dffeas \D_iw[29] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[29] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[29]~q ),
	.prn(vcc));
defparam \D_iw[29] .is_wysiwyg = "true";
defparam \D_iw[29] .power_up = "low";

dffeas \D_iw[31] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[31] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[31]~q ),
	.prn(vcc));
defparam \D_iw[31] .is_wysiwyg = "true";
defparam \D_iw[31] .power_up = "low";

dffeas \D_iw[30] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[30] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[30]~q ),
	.prn(vcc));
defparam \D_iw[30] .is_wysiwyg = "true";
defparam \D_iw[30] .power_up = "low";

dffeas \D_iw[27] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[27] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\F_iw~0_combout ),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[27]~q ),
	.prn(vcc));
defparam \D_iw[27] .is_wysiwyg = "true";
defparam \D_iw[27] .power_up = "low";

cyclonev_lcell_comb \Equal296~0 (
	.dataa(!\D_iw[28]~q ),
	.datab(!\D_iw[29]~q ),
	.datac(!\D_iw[31]~q ),
	.datad(!\D_iw[30]~q ),
	.datae(!\D_iw[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal296~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal296~0 .extended_lut = "off";
defparam \Equal296~0 .lut_mask = 64'hFFFFFFFEFFFFFFFE;
defparam \Equal296~0 .shared_arith = "off";

cyclonev_lcell_comb D_src1_hazard_E(
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\E_regnum_a_cmp_D~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_hazard_E~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_src1_hazard_E.extended_lut = "off";
defparam D_src1_hazard_E.lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam D_src1_hazard_E.shared_arith = "off";

dffeas \E_src1[4] (
	.clk(clk_clk),
	.d(\D_src1_reg[4]~10_combout ),
	.asdata(\E_alu_result[4]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[4]~q ),
	.prn(vcc));
defparam \E_src1[4] .is_wysiwyg = "true";
defparam \E_src1[4] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[1]~30 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[1] ),
	.datab(!\W_wr_data[1]~q ),
	.datac(!\M_alu_result[1]~q ),
	.datad(!\A_wr_data_unfiltered[1]~29_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[1]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[1]~30 .extended_lut = "off";
defparam \D_src1_reg[1]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[1]~30 .shared_arith = "off";

dffeas \E_src1[1] (
	.clk(clk_clk),
	.d(\D_src1_reg[1]~30_combout ),
	.asdata(\E_alu_result[1]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[1]~q ),
	.prn(vcc));
defparam \E_src1[1] .is_wysiwyg = "true";
defparam \E_src1[1] .power_up = "low";

dffeas \d_readdata_d1[0] (
	.clk(clk_clk),
	.d(d_readdata[0]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[0]~q ),
	.prn(vcc));
defparam \d_readdata_d1[0] .is_wysiwyg = "true";
defparam \d_readdata_d1[0] .power_up = "low";

dffeas \d_readdata_d1[8] (
	.clk(clk_clk),
	.d(d_readdata[8]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[8]~q ),
	.prn(vcc));
defparam \d_readdata_d1[8] .is_wysiwyg = "true";
defparam \d_readdata_d1[8] .power_up = "low";

dffeas \d_readdata_d1[16] (
	.clk(clk_clk),
	.d(d_readdata[16]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[16]~q ),
	.prn(vcc));
defparam \d_readdata_d1[16] .is_wysiwyg = "true";
defparam \d_readdata_d1[16] .power_up = "low";

dffeas \d_readdata_d1[24] (
	.clk(clk_clk),
	.d(d_readdata[24]),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\d_readdata_d1[24]~q ),
	.prn(vcc));
defparam \d_readdata_d1[24] .is_wysiwyg = "true";
defparam \d_readdata_d1[24] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte0_data_aligned_nxt[0]~7 (
	.dataa(!\d_readdata_d1[0]~q ),
	.datab(!\d_readdata_d1[8]~q ),
	.datac(!\d_readdata_d1[16]~q ),
	.datad(!\d_readdata_d1[24]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte0_data_aligned_nxt[0]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte0_data_aligned_nxt[0]~7 .extended_lut = "off";
defparam \A_slow_ld_byte0_data_aligned_nxt[0]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_ld_byte0_data_aligned_nxt[0]~7 .shared_arith = "off";

dffeas \A_slow_inst_result[0] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte0_data_aligned_nxt[0]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[0]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[0] .is_wysiwyg = "true";
defparam \A_slow_inst_result[0] .power_up = "low";

cyclonev_lcell_comb \M_inst_result~0 (
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\M_ctrl_mem~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[0] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_inst_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_inst_result~0 .extended_lut = "off";
defparam \M_inst_result~0 .lut_mask = 64'h4747474747474747;
defparam \M_inst_result~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_crst~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[15]~q ),
	.datae(!\D_ctrl_logic~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_crst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_crst~0 .extended_lut = "off";
defparam \D_ctrl_crst~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \D_ctrl_crst~0 .shared_arith = "off";

dffeas E_ctrl_crst(
	.clk(clk_clk),
	.d(\D_ctrl_crst~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_crst~q ),
	.prn(vcc));
defparam E_ctrl_crst.is_wysiwyg = "true";
defparam E_ctrl_crst.power_up = "low";

dffeas M_ctrl_crst(
	.clk(clk_clk),
	.d(\E_ctrl_crst~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_crst~q ),
	.prn(vcc));
defparam M_ctrl_crst.is_wysiwyg = "true";
defparam M_ctrl_crst.power_up = "low";

cyclonev_lcell_comb \D_ctrl_break~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[15]~q ),
	.datae(!\D_ctrl_logic~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_break~0 .extended_lut = "off";
defparam \D_ctrl_break~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \D_ctrl_break~0 .shared_arith = "off";

dffeas E_ctrl_break(
	.clk(clk_clk),
	.d(\D_ctrl_break~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_break~q ),
	.prn(vcc));
defparam E_ctrl_break.is_wysiwyg = "true";
defparam E_ctrl_break.power_up = "low";

dffeas M_ctrl_break(
	.clk(clk_clk),
	.d(\E_ctrl_break~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_break~q ),
	.prn(vcc));
defparam M_ctrl_break.is_wysiwyg = "true";
defparam M_ctrl_break.power_up = "low";

cyclonev_lcell_comb \D_ctrl_exception~0 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[11]~q ),
	.datad(!\D_iw[16]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_ctrl_logic~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_exception~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_exception~0 .extended_lut = "off";
defparam \D_ctrl_exception~0 .lut_mask = 64'h6F9F9F6FFFFFFFFF;
defparam \D_ctrl_exception~0 .shared_arith = "off";

dffeas E_ctrl_exception(
	.clk(clk_clk),
	.d(\D_ctrl_exception~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_exception~q ),
	.prn(vcc));
defparam E_ctrl_exception.is_wysiwyg = "true";
defparam E_ctrl_exception.power_up = "low";

dffeas M_ctrl_exception(
	.clk(clk_clk),
	.d(\E_ctrl_exception~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_exception~q ),
	.prn(vcc));
defparam M_ctrl_exception.is_wysiwyg = "true";
defparam M_ctrl_exception.power_up = "low";

dffeas \M_iw[14] (
	.clk(clk_clk),
	.d(\E_iw[14]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[14]~q ),
	.prn(vcc));
defparam \M_iw[14] .is_wysiwyg = "true";
defparam \M_iw[14] .power_up = "low";

dffeas \M_iw[11] (
	.clk(clk_clk),
	.d(\E_iw[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[11]~q ),
	.prn(vcc));
defparam \M_iw[11] .is_wysiwyg = "true";
defparam \M_iw[11] .power_up = "low";

dffeas \M_iw[5] (
	.clk(clk_clk),
	.d(\E_iw[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[5]~q ),
	.prn(vcc));
defparam \M_iw[5] .is_wysiwyg = "true";
defparam \M_iw[5] .power_up = "low";

dffeas \M_iw[0] (
	.clk(clk_clk),
	.d(\E_iw[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[0]~q ),
	.prn(vcc));
defparam \M_iw[0] .is_wysiwyg = "true";
defparam \M_iw[0] .power_up = "low";

dffeas \M_iw[16] (
	.clk(clk_clk),
	.d(\E_iw[16]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[16]~q ),
	.prn(vcc));
defparam \M_iw[16] .is_wysiwyg = "true";
defparam \M_iw[16] .power_up = "low";

dffeas \M_iw[15] (
	.clk(clk_clk),
	.d(\E_iw[15]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[15]~q ),
	.prn(vcc));
defparam \M_iw[15] .is_wysiwyg = "true";
defparam \M_iw[15] .power_up = "low";

dffeas \M_iw[13] (
	.clk(clk_clk),
	.d(\E_iw[13]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[13]~q ),
	.prn(vcc));
defparam \M_iw[13] .is_wysiwyg = "true";
defparam \M_iw[13] .power_up = "low";

dffeas \M_iw[12] (
	.clk(clk_clk),
	.d(\E_iw[12]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[12]~q ),
	.prn(vcc));
defparam \M_iw[12] .is_wysiwyg = "true";
defparam \M_iw[12] .power_up = "low";

cyclonev_lcell_comb \M_op_eret~0 (
	.dataa(!\M_iw[16]~q ),
	.datab(!\M_iw[15]~q ),
	.datac(!\M_iw[13]~q ),
	.datad(!\M_iw[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_op_eret~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_op_eret~0 .extended_lut = "off";
defparam \M_op_eret~0 .lut_mask = 64'hFFFEFFFEFFFEFFFE;
defparam \M_op_eret~0 .shared_arith = "off";

dffeas \M_iw[4] (
	.clk(clk_clk),
	.d(\E_iw[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[4]~q ),
	.prn(vcc));
defparam \M_iw[4] .is_wysiwyg = "true";
defparam \M_iw[4] .power_up = "low";

dffeas \M_iw[3] (
	.clk(clk_clk),
	.d(\E_iw[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[3]~q ),
	.prn(vcc));
defparam \M_iw[3] .is_wysiwyg = "true";
defparam \M_iw[3] .power_up = "low";

dffeas \M_iw[2] (
	.clk(clk_clk),
	.d(\E_iw[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[2]~q ),
	.prn(vcc));
defparam \M_iw[2] .is_wysiwyg = "true";
defparam \M_iw[2] .power_up = "low";

dffeas \M_iw[1] (
	.clk(clk_clk),
	.d(\E_iw[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[1]~q ),
	.prn(vcc));
defparam \M_iw[1] .is_wysiwyg = "true";
defparam \M_iw[1] .power_up = "low";

cyclonev_lcell_comb \M_op_eret~1 (
	.dataa(!\M_iw[4]~q ),
	.datab(!\M_iw[3]~q ),
	.datac(!\M_iw[2]~q ),
	.datad(!\M_iw[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_op_eret~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_op_eret~1 .extended_lut = "off";
defparam \M_op_eret~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \M_op_eret~1 .shared_arith = "off";

cyclonev_lcell_comb \M_op_eret~2 (
	.dataa(!\M_iw[11]~q ),
	.datab(!\M_iw[5]~q ),
	.datac(!\M_iw[0]~q ),
	.datad(!\M_op_eret~0_combout ),
	.datae(!\M_op_eret~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_op_eret~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_op_eret~2 .extended_lut = "off";
defparam \M_op_eret~2 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \M_op_eret~2 .shared_arith = "off";

dffeas \E_iw[6] (
	.clk(clk_clk),
	.d(\D_iw[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[6]~q ),
	.prn(vcc));
defparam \E_iw[6] .is_wysiwyg = "true";
defparam \E_iw[6] .power_up = "low";

dffeas \M_iw[6] (
	.clk(clk_clk),
	.d(\E_iw[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[6]~q ),
	.prn(vcc));
defparam \M_iw[6] .is_wysiwyg = "true";
defparam \M_iw[6] .power_up = "low";

dffeas \E_iw[7] (
	.clk(clk_clk),
	.d(\D_iw[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[7]~q ),
	.prn(vcc));
defparam \E_iw[7] .is_wysiwyg = "true";
defparam \E_iw[7] .power_up = "low";

dffeas \M_iw[7] (
	.clk(clk_clk),
	.d(\E_iw[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[7]~q ),
	.prn(vcc));
defparam \M_iw[7] .is_wysiwyg = "true";
defparam \M_iw[7] .power_up = "low";

dffeas \E_iw[8] (
	.clk(clk_clk),
	.d(\D_iw[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[8]~q ),
	.prn(vcc));
defparam \E_iw[8] .is_wysiwyg = "true";
defparam \E_iw[8] .power_up = "low";

dffeas \M_iw[8] (
	.clk(clk_clk),
	.d(\E_iw[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_iw[8]~q ),
	.prn(vcc));
defparam \M_iw[8] .is_wysiwyg = "true";
defparam \M_iw[8] .power_up = "low";

cyclonev_lcell_comb E_op_wrctl(
	.dataa(!\E_iw[14]~q ),
	.datab(!\E_op_rdctl~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_op_wrctl~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_op_wrctl.extended_lut = "off";
defparam E_op_wrctl.lut_mask = 64'h7777777777777777;
defparam E_op_wrctl.shared_arith = "off";

dffeas M_ctrl_wrctl_inst(
	.clk(clk_clk),
	.d(\E_op_wrctl~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_wrctl_inst~q ),
	.prn(vcc));
defparam M_ctrl_wrctl_inst.is_wysiwyg = "true";
defparam M_ctrl_wrctl_inst.power_up = "low";

cyclonev_lcell_comb M_wrctl_bstatus(
	.dataa(!\M_iw[6]~q ),
	.datab(!\M_iw[7]~q ),
	.datac(!\M_iw[8]~q ),
	.datad(!\M_ctrl_wrctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wrctl_bstatus~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_wrctl_bstatus.extended_lut = "off";
defparam M_wrctl_bstatus.lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam M_wrctl_bstatus.shared_arith = "off";

cyclonev_lcell_comb \A_bstatus_reg_pie_inst_nxt~0 (
	.dataa(!\M_ctrl_break~q ),
	.datab(!\M_alu_result[0]~q ),
	.datac(!\A_bstatus_reg_pie~q ),
	.datad(!\A_status_reg_pie~q ),
	.datae(!\M_wrctl_bstatus~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_bstatus_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_bstatus_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \A_bstatus_reg_pie_inst_nxt~0 .lut_mask = 64'h7FFFBFFF7FFFBFFF;
defparam \A_bstatus_reg_pie_inst_nxt~0 .shared_arith = "off";

dffeas A_bstatus_reg_pie(
	.clk(clk_clk),
	.d(\A_bstatus_reg_pie_inst_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always120~0_combout ),
	.q(\A_bstatus_reg_pie~q ),
	.prn(vcc));
defparam A_bstatus_reg_pie.is_wysiwyg = "true";
defparam A_bstatus_reg_pie.power_up = "low";

cyclonev_lcell_comb \A_status_reg_pie_inst_nxt~0 (
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\A_status_reg_pie~q ),
	.datac(!\M_iw[6]~q ),
	.datad(!\M_iw[7]~q ),
	.datae(!\M_iw[8]~q ),
	.dataf(!\M_ctrl_wrctl_inst~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_status_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_status_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \A_status_reg_pie_inst_nxt~0 .lut_mask = 64'h7FF7F77FF77F7FF7;
defparam \A_status_reg_pie_inst_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \A_status_reg_pie_inst_nxt~1 (
	.dataa(!\M_iw[14]~q ),
	.datab(!\M_op_eret~2_combout ),
	.datac(!\A_estatus_reg_pie~q ),
	.datad(!\A_bstatus_reg_pie~q ),
	.datae(!\A_status_reg_pie_inst_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_status_reg_pie_inst_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_status_reg_pie_inst_nxt~1 .extended_lut = "off";
defparam \A_status_reg_pie_inst_nxt~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_status_reg_pie_inst_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \A_status_reg_pie_inst_nxt~2 (
	.dataa(!\M_ctrl_break~q ),
	.datab(!\M_ctrl_crst~q ),
	.datac(!\M_ctrl_exception~q ),
	.datad(!\A_status_reg_pie_inst_nxt~1_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_status_reg_pie_inst_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_status_reg_pie_inst_nxt~2 .extended_lut = "off";
defparam \A_status_reg_pie_inst_nxt~2 .lut_mask = 64'hFEFFFEFFFEFFFEFF;
defparam \A_status_reg_pie_inst_nxt~2 .shared_arith = "off";

dffeas A_status_reg_pie(
	.clk(clk_clk),
	.d(\A_status_reg_pie_inst_nxt~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always120~0_combout ),
	.q(\A_status_reg_pie~q ),
	.prn(vcc));
defparam A_status_reg_pie.is_wysiwyg = "true";
defparam A_status_reg_pie.power_up = "low";

cyclonev_lcell_comb M_wrctl_estatus(
	.dataa(!\M_iw[6]~q ),
	.datab(!\M_iw[7]~q ),
	.datac(!\M_iw[8]~q ),
	.datad(!\M_ctrl_wrctl_inst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_wrctl_estatus~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_wrctl_estatus.extended_lut = "off";
defparam M_wrctl_estatus.lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam M_wrctl_estatus.shared_arith = "off";

cyclonev_lcell_comb \A_estatus_reg_pie_inst_nxt~0 (
	.dataa(!\M_alu_result[0]~q ),
	.datab(!\M_ctrl_crst~q ),
	.datac(!\A_estatus_reg_pie~q ),
	.datad(!\A_status_reg_pie~q ),
	.datae(!\M_ctrl_exception~q ),
	.dataf(!\M_wrctl_estatus~combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_estatus_reg_pie_inst_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_estatus_reg_pie_inst_nxt~0 .extended_lut = "off";
defparam \A_estatus_reg_pie_inst_nxt~0 .lut_mask = 64'hDFFFFFFFFFFFDFFF;
defparam \A_estatus_reg_pie_inst_nxt~0 .shared_arith = "off";

dffeas A_estatus_reg_pie(
	.clk(clk_clk),
	.d(\A_estatus_reg_pie_inst_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always120~0_combout ),
	.q(\A_estatus_reg_pie~q ),
	.prn(vcc));
defparam A_estatus_reg_pie.is_wysiwyg = "true";
defparam A_estatus_reg_pie.power_up = "low";

cyclonev_lcell_comb \D_control_reg_rddata_muxed[0]~0 (
	.dataa(!\D_iw[8]~q ),
	.datab(!\D_iw[6]~q ),
	.datac(!\D_iw[7]~q ),
	.datad(!\A_estatus_reg_pie~q ),
	.datae(!\A_bstatus_reg_pie~q ),
	.dataf(!\A_status_reg_pie~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_control_reg_rddata_muxed[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_control_reg_rddata_muxed[0]~0 .extended_lut = "off";
defparam \D_control_reg_rddata_muxed[0]~0 .lut_mask = 64'hBEFFFFFFFFFFFFFF;
defparam \D_control_reg_rddata_muxed[0]~0 .shared_arith = "off";

dffeas \E_control_reg_rddata[0] (
	.clk(clk_clk),
	.d(\D_control_reg_rddata_muxed[0]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_control_reg_rddata[0]~q ),
	.prn(vcc));
defparam \E_control_reg_rddata[0] .is_wysiwyg = "true";
defparam \E_control_reg_rddata[0] .power_up = "low";

dffeas \M_control_reg_rddata[0] (
	.clk(clk_clk),
	.d(\E_control_reg_rddata[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_control_reg_rddata[0]~q ),
	.prn(vcc));
defparam \M_control_reg_rddata[0] .is_wysiwyg = "true";
defparam \M_control_reg_rddata[0] .power_up = "low";

dffeas \A_inst_result[0] (
	.clk(clk_clk),
	.d(\M_inst_result~0_combout ),
	.asdata(\M_control_reg_rddata[0]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\M_ctrl_rdctl_inst~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[0]~q ),
	.prn(vcc));
defparam \A_inst_result[0] .is_wysiwyg = "true";
defparam \A_inst_result[0] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[0]~5 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[0]~5 .extended_lut = "off";
defparam \E_rot_mask[0]~5 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[0]~5 .shared_arith = "off";

dffeas \M_rot_mask[0] (
	.clk(clk_clk),
	.d(\E_rot_mask[0]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[0]~q ),
	.prn(vcc));
defparam \M_rot_mask[0] .is_wysiwyg = "true";
defparam \M_rot_mask[0] .power_up = "low";

cyclonev_lcell_comb \Add7~0 (
	.dataa(!\E_src2[1]~q ),
	.datab(!\E_src2[0]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~0 .extended_lut = "off";
defparam \Add7~0 .lut_mask = 64'h9696969696969696;
defparam \Add7~0 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[4]~19 (
	.dataa(!\E_src1[4]~q ),
	.datab(!\E_src1[3]~q ),
	.datac(!\E_src1[2]~q ),
	.datad(!\E_src1[1]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[4]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[4]~19 .extended_lut = "off";
defparam \E_rot_step1[4]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[4]~19 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_reg[8]~6 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[8] ),
	.datab(!\W_wr_data[8]~q ),
	.datac(!\M_alu_result[8]~q ),
	.datad(!\A_wr_data_unfiltered[8]~17_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[8]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[8]~6 .extended_lut = "off";
defparam \D_src1_reg[8]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[8]~6 .shared_arith = "off";

dffeas \E_src1[8] (
	.clk(clk_clk),
	.d(\D_src1_reg[8]~6_combout ),
	.asdata(\E_alu_result[8]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[8]~q ),
	.prn(vcc));
defparam \E_src1[8] .is_wysiwyg = "true";
defparam \E_src1[8] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[8]~16 (
	.dataa(!\E_src1[8]~q ),
	.datab(!\E_src1[7]~q ),
	.datac(!\E_src1[6]~q ),
	.datad(!\E_src1[5]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[8]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[8]~16 .extended_lut = "off";
defparam \E_rot_step1[8]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[8]~16 .shared_arith = "off";

cyclonev_lcell_comb \Add7~1 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~1 .extended_lut = "off";
defparam \Add7~1 .lut_mask = 64'h6996699669966996;
defparam \Add7~1 .shared_arith = "off";

dffeas \M_rot_prestep2[8] (
	.clk(clk_clk),
	.d(\E_rot_step1[4]~19_combout ),
	.asdata(\E_rot_step1[8]~16_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[8]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[8] .is_wysiwyg = "true";
defparam \M_rot_prestep2[8] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[17]~16 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[17] ),
	.datab(!\W_wr_data[17]~q ),
	.datac(!\M_alu_result[17]~q ),
	.datad(!\A_wr_data_unfiltered[17]~40_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[17]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[17]~16 .extended_lut = "off";
defparam \D_src1_reg[17]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[17]~16 .shared_arith = "off";

dffeas \E_src1[17] (
	.clk(clk_clk),
	.d(\D_src1_reg[17]~16_combout ),
	.asdata(\E_alu_result[17]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[17]~q ),
	.prn(vcc));
defparam \E_src1[17] .is_wysiwyg = "true";
defparam \E_src1[17] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~17 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[17]~q ),
	.datae(!\E_src1[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~17 .extended_lut = "off";
defparam \E_alu_result~17 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~17 .shared_arith = "off";

cyclonev_lcell_comb \D_src1_reg[16]~17 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[16] ),
	.datab(!\W_wr_data[16]~q ),
	.datac(!\M_alu_result[16]~q ),
	.datad(!\A_wr_data_unfiltered[16]~44_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[16]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[16]~17 .extended_lut = "off";
defparam \D_src1_reg[16]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[16]~17 .shared_arith = "off";

dffeas \E_src1[16] (
	.clk(clk_clk),
	.d(\D_src1_reg[16]~17_combout ),
	.asdata(\E_alu_result[16]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[16]~q ),
	.prn(vcc));
defparam \E_src1[16] .is_wysiwyg = "true";
defparam \E_src1[16] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~19 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[16]~q ),
	.datae(!\E_src1[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~19 .extended_lut = "off";
defparam \E_alu_result~19 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~19 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_mask[7]~6 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[7]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[7]~6 .extended_lut = "off";
defparam \E_rot_mask[7]~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[7]~6 .shared_arith = "off";

dffeas \M_rot_mask[7] (
	.clk(clk_clk),
	.d(\E_rot_mask[7]~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[7]~q ),
	.prn(vcc));
defparam \M_rot_mask[7] .is_wysiwyg = "true";
defparam \M_rot_mask[7] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[11]~3 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[11] ),
	.datab(!\W_wr_data[11]~q ),
	.datac(!\M_alu_result[11]~q ),
	.datad(!\A_wr_data_unfiltered[11]~11_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[11]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[11]~3 .extended_lut = "off";
defparam \D_src1_reg[11]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[11]~3 .shared_arith = "off";

dffeas \E_src1[11] (
	.clk(clk_clk),
	.d(\D_src1_reg[11]~3_combout ),
	.asdata(\E_alu_result[11]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[11]~q ),
	.prn(vcc));
defparam \E_src1[11] .is_wysiwyg = "true";
defparam \E_src1[11] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[1]~4 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[1]~4 .extended_lut = "off";
defparam \E_rot_mask[1]~4 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[1]~4 .shared_arith = "off";

dffeas \M_rot_mask[1] (
	.clk(clk_clk),
	.d(\E_rot_mask[1]~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[1]~q ),
	.prn(vcc));
defparam \M_rot_mask[1] .is_wysiwyg = "true";
defparam \M_rot_mask[1] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[5]~11 (
	.dataa(!\E_src1[5]~q ),
	.datab(!\E_src1[4]~q ),
	.datac(!\E_src1[3]~q ),
	.datad(!\E_src1[2]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[5]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[5]~11 .extended_lut = "off";
defparam \E_rot_step1[5]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[5]~11 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[9]~8 (
	.dataa(!\E_src1[9]~q ),
	.datab(!\E_src1[8]~q ),
	.datac(!\E_src1[7]~q ),
	.datad(!\E_src1[6]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[9]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[9]~8 .extended_lut = "off";
defparam \E_rot_step1[9]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[9]~8 .shared_arith = "off";

dffeas \M_rot_prestep2[9] (
	.clk(clk_clk),
	.d(\E_rot_step1[5]~11_combout ),
	.asdata(\E_rot_step1[9]~8_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[9]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[9] .is_wysiwyg = "true";
defparam \M_rot_prestep2[9] .power_up = "low";

cyclonev_lcell_comb \Add17~133 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[28]~q ),
	.datae(gnd),
	.dataf(!\E_src1[28]~q ),
	.datag(gnd),
	.cin(\Add17~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~133_sumout ),
	.cout(\Add17~134 ),
	.shareout());
defparam \Add17~133 .extended_lut = "off";
defparam \Add17~133 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~133 .shared_arith = "off";

cyclonev_lcell_comb \Add17~129 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[29]~q ),
	.datae(gnd),
	.dataf(!\E_src1[29]~q ),
	.datag(gnd),
	.cin(\Add17~134 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~129_sumout ),
	.cout(\Add17~130 ),
	.shareout());
defparam \Add17~129 .extended_lut = "off";
defparam \Add17~129 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~129 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~57 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~28_combout ),
	.datad(!\Add17~129_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~57 .extended_lut = "off";
defparam \D_src2_reg[29]~57 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[29]~57 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~58 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[29]~q ),
	.datae(!\A_wr_data_unfiltered[29]~60_combout ),
	.dataf(!\M_alu_result[29]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~58 .extended_lut = "off";
defparam \D_src2_reg[29]~58 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[29]~58 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_unsigned_lo_imm16~1 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[1] ),
	.datac(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[5] ),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[3] ),
	.datae(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[2] ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_unsigned_lo_imm16~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_unsigned_lo_imm16~1 .extended_lut = "off";
defparam \F_ctrl_unsigned_lo_imm16~1 .lut_mask = 64'hEFFEFEEFFEEFEFFE;
defparam \F_ctrl_unsigned_lo_imm16~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ctrl_unsigned_lo_imm16~0 (
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[12]~11_combout ),
	.datac(!\F_iw[11]~12_combout ),
	.datad(!\F_iw[13]~8_combout ),
	.datae(!\Equal2~0_combout ),
	.dataf(!\F_ctrl_unsigned_lo_imm16~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_unsigned_lo_imm16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_unsigned_lo_imm16~0 .extended_lut = "off";
defparam \F_ctrl_unsigned_lo_imm16~0 .lut_mask = 64'hFFFBFFFFFFFFFFFF;
defparam \F_ctrl_unsigned_lo_imm16~0 .shared_arith = "off";

dffeas D_ctrl_unsigned_lo_imm16(
	.clk(clk_clk),
	.d(\F_ctrl_unsigned_lo_imm16~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_unsigned_lo_imm16~q ),
	.prn(vcc));
defparam D_ctrl_unsigned_lo_imm16.is_wysiwyg = "true";
defparam D_ctrl_unsigned_lo_imm16.power_up = "low";

cyclonev_lcell_comb \D_src2[29]~2 (
	.dataa(!\D_iw[19]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[29]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[29]~2 .extended_lut = "off";
defparam \D_src2[29]~2 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[29]~2 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[29]~3 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[29]~57_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.datae(!\D_src2_reg[29]~58_combout ),
	.dataf(!\D_src2[29]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[29]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[29]~3 .extended_lut = "off";
defparam \D_src2[29]~3 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[29]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_src2[19]~1 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_src2[19]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_src2[19]~1 .extended_lut = "off";
defparam \E_src2[19]~1 .lut_mask = 64'h7777777777777777;
defparam \E_src2[19]~1 .shared_arith = "off";

dffeas \E_src2[29] (
	.clk(clk_clk),
	.d(\D_src2[29]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[29]~q ),
	.prn(vcc));
defparam \E_src2[29] .is_wysiwyg = "true";
defparam \E_src2[29] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[29]~7 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[29]~q ),
	.datad(!\E_src1[29]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[29]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[29]~7 .extended_lut = "off";
defparam \E_logic_result[29]~7 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[29]~7 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~28 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[29]~7_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~28 .extended_lut = "off";
defparam \E_alu_result~28 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~28 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[29] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~28_combout ),
	.datac(!\Add17~129_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[29]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[29] .extended_lut = "off";
defparam \E_alu_result[29] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[29] .shared_arith = "off";

dffeas \M_alu_result[29] (
	.clk(clk_clk),
	.d(\E_alu_result[29]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[29]~q ),
	.prn(vcc));
defparam \M_alu_result[29] .is_wysiwyg = "true";
defparam \M_alu_result[29] .power_up = "low";

dffeas \A_inst_result[29] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[29] ),
	.asdata(\M_alu_result[29]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[29]~q ),
	.prn(vcc));
defparam \A_inst_result[29] .is_wysiwyg = "true";
defparam \A_inst_result[29] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[5]~1 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[5]~1 .extended_lut = "off";
defparam \E_rot_mask[5]~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[5]~1 .shared_arith = "off";

dffeas \M_rot_mask[5] (
	.clk(clk_clk),
	.d(\E_rot_mask[5]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[5]~q ),
	.prn(vcc));
defparam \M_rot_mask[5] .is_wysiwyg = "true";
defparam \M_rot_mask[5] .power_up = "low";

cyclonev_lcell_comb \D_ctrl_rot~0 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\Equal171~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_rot~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_rot~0 .extended_lut = "off";
defparam \D_ctrl_rot~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \D_ctrl_rot~0 .shared_arith = "off";

dffeas E_ctrl_rot(
	.clk(clk_clk),
	.d(\D_ctrl_rot~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_rot~q ),
	.prn(vcc));
defparam E_ctrl_rot.is_wysiwyg = "true";
defparam E_ctrl_rot.power_up = "low";

cyclonev_lcell_comb \E_rot_pass3~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_left~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass3~0 .extended_lut = "off";
defparam \E_rot_pass3~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \E_rot_pass3~0 .shared_arith = "off";

dffeas M_rot_pass3(
	.clk(clk_clk),
	.d(\E_rot_pass3~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_pass3~q ),
	.prn(vcc));
defparam M_rot_pass3.is_wysiwyg = "true";
defparam M_rot_pass3.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill3~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill3~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill3~0 .extended_lut = "off";
defparam \E_rot_sel_fill3~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_rot_sel_fill3~0 .shared_arith = "off";

dffeas M_rot_sel_fill3(
	.clk(clk_clk),
	.d(\E_rot_sel_fill3~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_sel_fill3~q ),
	.prn(vcc));
defparam M_rot_sel_fill3.is_wysiwyg = "true";
defparam M_rot_sel_fill3.power_up = "low";

cyclonev_lcell_comb \E_rot_step1[25]~12 (
	.dataa(!\E_src1[25]~q ),
	.datab(!\E_src1[24]~q ),
	.datac(!\E_src1[23]~q ),
	.datad(!\E_src1[22]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[25]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[25]~12 .extended_lut = "off";
defparam \E_rot_step1[25]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[25]~12 .shared_arith = "off";

dffeas \M_rot_prestep2[29] (
	.clk(clk_clk),
	.d(\E_rot_step1[25]~12_combout ),
	.asdata(\E_rot_step1[29]~13_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[29]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[29] .is_wysiwyg = "true";
defparam \M_rot_prestep2[29] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[14]~27 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[14] ),
	.datab(!\W_wr_data[14]~q ),
	.datac(!\M_alu_result[14]~q ),
	.datad(!\A_wr_data_unfiltered[14]~68_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[14]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[14]~27 .extended_lut = "off";
defparam \D_src1_reg[14]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[14]~27 .shared_arith = "off";

dffeas \E_src1[14] (
	.clk(clk_clk),
	.d(\D_src1_reg[14]~27_combout ),
	.asdata(\E_alu_result[14]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[14]~q ),
	.prn(vcc));
defparam \E_src1[14] .is_wysiwyg = "true";
defparam \E_src1[14] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[17]~14 (
	.dataa(!\E_src1[17]~q ),
	.datab(!\E_src1[16]~q ),
	.datac(!\E_src1[15]~q ),
	.datad(!\E_src1[14]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[17]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[17]~14 .extended_lut = "off";
defparam \E_rot_step1[17]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[17]~14 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[21]~15 (
	.dataa(!\E_src1[21]~q ),
	.datab(!\E_src1[20]~q ),
	.datac(!\E_src1[19]~q ),
	.datad(!\E_src1[18]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[21]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[21]~15 .extended_lut = "off";
defparam \E_rot_step1[21]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[21]~15 .shared_arith = "off";

dffeas \M_rot_prestep2[21] (
	.clk(clk_clk),
	.d(\E_rot_step1[17]~14_combout ),
	.asdata(\E_rot_step1[21]~15_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[21]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[21] .is_wysiwyg = "true";
defparam \M_rot_prestep2[21] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[30]~8 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[30]~q ),
	.datad(!\E_src1[30]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[30]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[30]~8 .extended_lut = "off";
defparam \E_logic_result[30]~8 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[30]~8 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~29 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[30]~8_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~29 .extended_lut = "off";
defparam \E_alu_result~29 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~29 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[30]~59 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add17~65_sumout ),
	.datac(!\D_src2_reg[0]~28_combout ),
	.datad(!\E_alu_result~29_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~59 .extended_lut = "off";
defparam \D_src2_reg[30]~59 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[30]~59 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[30]~60 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[30]~q ),
	.datae(!\A_wr_data_unfiltered[30]~62_combout ),
	.dataf(!\M_alu_result[30]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~60 .extended_lut = "off";
defparam \D_src2_reg[30]~60 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[30]~60 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[30]~4 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[21]~q ),
	.datac(!\D_iw[20]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[30]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[30]~4 .extended_lut = "off";
defparam \D_src2[30]~4 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \D_src2[30]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[30]~5 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[30]~59_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.datae(!\D_src2_reg[30]~60_combout ),
	.dataf(!\D_src2[30]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[30]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[30]~5 .extended_lut = "off";
defparam \D_src2[30]~5 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[30]~5 .shared_arith = "off";

dffeas \E_src2[30] (
	.clk(clk_clk),
	.d(\D_src2[30]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[30]~q ),
	.prn(vcc));
defparam \E_src2[30] .is_wysiwyg = "true";
defparam \E_src2[30] .power_up = "low";

cyclonev_lcell_comb \Add17~65 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[30]~q ),
	.datae(gnd),
	.dataf(!\E_src1[30]~q ),
	.datag(gnd),
	.cin(\Add17~130 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~65_sumout ),
	.cout(\Add17~66 ),
	.shareout());
defparam \Add17~65 .extended_lut = "off";
defparam \Add17~65 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~65 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[30] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add17~65_sumout ),
	.datac(!\E_alu_result~29_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[30]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[30] .extended_lut = "off";
defparam \E_alu_result[30] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[30] .shared_arith = "off";

dffeas \M_alu_result[30] (
	.clk(clk_clk),
	.d(\E_alu_result[30]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[30]~q ),
	.prn(vcc));
defparam \M_alu_result[30] .is_wysiwyg = "true";
defparam \M_alu_result[30] .power_up = "low";

dffeas \A_inst_result[30] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[30] ),
	.asdata(\M_alu_result[30]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[30]~q ),
	.prn(vcc));
defparam \A_inst_result[30] .is_wysiwyg = "true";
defparam \A_inst_result[30] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[26]~3 (
	.dataa(!\E_src1[26]~q ),
	.datab(!\E_src1[25]~q ),
	.datac(!\E_src1[24]~q ),
	.datad(!\E_src1[23]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[26]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[26]~3 .extended_lut = "off";
defparam \E_rot_step1[26]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[26]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[30]~0 (
	.dataa(!\E_src1[30]~q ),
	.datab(!\E_src1[29]~q ),
	.datac(!\E_src1[28]~q ),
	.datad(!\E_src1[27]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[30]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[30]~0 .extended_lut = "off";
defparam \E_rot_step1[30]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[30]~0 .shared_arith = "off";

dffeas \M_rot_prestep2[30] (
	.clk(clk_clk),
	.d(\E_rot_step1[26]~3_combout ),
	.asdata(\E_rot_step1[30]~0_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[30]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[30] .is_wysiwyg = "true";
defparam \M_rot_prestep2[30] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[18]~5 (
	.dataa(!\E_src1[18]~q ),
	.datab(!\E_src1[17]~q ),
	.datac(!\E_src1[16]~q ),
	.datad(!\E_src1[15]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[18]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[18]~5 .extended_lut = "off";
defparam \E_rot_step1[18]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[18]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[22]~2 (
	.dataa(!\E_src1[22]~q ),
	.datab(!\E_src1[21]~q ),
	.datac(!\E_src1[20]~q ),
	.datad(!\E_src1[19]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[22]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[22]~2 .extended_lut = "off";
defparam \E_rot_step1[22]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[22]~2 .shared_arith = "off";

dffeas \M_rot_prestep2[22] (
	.clk(clk_clk),
	.d(\E_rot_step1[18]~5_combout ),
	.asdata(\E_rot_step1[22]~2_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[22]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[22] .is_wysiwyg = "true";
defparam \M_rot_prestep2[22] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[2]~1 (
	.dataa(!\E_src1[2]~q ),
	.datab(!\E_src1[1]~q ),
	.datac(!\E_src1[0]~q ),
	.datad(!\E_src1[31]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[2]~1 .extended_lut = "off";
defparam \E_rot_step1[2]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[2]~1 .shared_arith = "off";

dffeas \M_rot_prestep2[6] (
	.clk(clk_clk),
	.d(\E_rot_step1[2]~1_combout ),
	.asdata(\E_rot_step1[6]~6_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[6]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[6] .is_wysiwyg = "true";
defparam \M_rot_prestep2[6] .power_up = "low";

cyclonev_lcell_comb \Add7~2 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_src2[3]~q ),
	.datae(!\E_ctrl_shift_rot_right~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~2 .extended_lut = "off";
defparam \Add7~2 .lut_mask = 64'h9669699696696996;
defparam \Add7~2 .shared_arith = "off";

dffeas \M_rot_rn[3] (
	.clk(clk_clk),
	.d(\Add7~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_rn[3]~q ),
	.prn(vcc));
defparam \M_rot_rn[3] .is_wysiwyg = "true";
defparam \M_rot_rn[3] .power_up = "low";

cyclonev_lcell_comb \Add7~3 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_src2[3]~q ),
	.datae(!\E_src2[4]~q ),
	.dataf(!\E_ctrl_shift_rot_right~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add7~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add7~3 .extended_lut = "off";
defparam \Add7~3 .lut_mask = 64'h6996966996696996;
defparam \Add7~3 .shared_arith = "off";

dffeas \M_rot_rn[4] (
	.clk(clk_clk),
	.d(\Add7~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_rn[4]~q ),
	.prn(vcc));
defparam \M_rot_rn[4] .is_wysiwyg = "true";
defparam \M_rot_rn[4] .power_up = "low";

cyclonev_lcell_comb \M_rot[6]~29 (
	.dataa(!\M_rot_prestep2[30]~q ),
	.datab(!\M_rot_prestep2[22]~q ),
	.datac(!\M_rot_prestep2[14]~q ),
	.datad(!\M_rot_prestep2[6]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~29 .extended_lut = "off";
defparam \M_rot[6]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~29 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~29 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[6]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[6]~29_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~29 .extended_lut = "off";
defparam \A_shift_rot_result~29 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~29 .shared_arith = "off";

dffeas \A_shift_rot_result[30] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~29_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[30]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[30] .is_wysiwyg = "true";
defparam \A_shift_rot_result[30] .power_up = "low";

dffeas \A_mem_baddr[1] (
	.clk(clk_clk),
	.d(\M_alu_result[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[1]~q ),
	.prn(vcc));
defparam \A_mem_baddr[1] .is_wysiwyg = "true";
defparam \A_mem_baddr[1] .power_up = "low";

dffeas \A_mem_baddr[0] (
	.clk(clk_clk),
	.d(\M_alu_result[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[0]~q ),
	.prn(vcc));
defparam \A_mem_baddr[0] .is_wysiwyg = "true";
defparam \A_mem_baddr[0] .power_up = "low";

cyclonev_lcell_comb \Equal187~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\E_iw[1]~q ),
	.datad(!\E_iw[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal187~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal187~0 .extended_lut = "off";
defparam \Equal187~0 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \Equal187~0 .shared_arith = "off";

dffeas M_ctrl_ld16(
	.clk(clk_clk),
	.d(\Equal187~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld16~q ),
	.prn(vcc));
defparam M_ctrl_ld16.is_wysiwyg = "true";
defparam M_ctrl_ld16.power_up = "low";

dffeas A_ctrl_ld16(
	.clk(clk_clk),
	.d(\M_ctrl_ld16~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_ld16~q ),
	.prn(vcc));
defparam A_ctrl_ld16.is_wysiwyg = "true";
defparam A_ctrl_ld16.power_up = "low";

cyclonev_lcell_comb \A_slow_ld_data_sign_bit~0 (
	.dataa(!\A_mem_baddr[0]~q ),
	.datab(!\A_ctrl_ld16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_data_sign_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_data_sign_bit~0 .extended_lut = "off";
defparam \A_slow_ld_data_sign_bit~0 .lut_mask = 64'h7777777777777777;
defparam \A_slow_ld_data_sign_bit~0 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_ld_data_fill_bit~0 (
	.dataa(!\A_mem_baddr[1]~q ),
	.datab(!\d_readdata_d1[31]~q ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\d_readdata_d1[23]~q ),
	.datae(!\A_slow_ld_data_sign_bit~0_combout ),
	.dataf(!\A_ctrl_ld_signed~q ),
	.datag(!\d_readdata_d1[7]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_data_fill_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_data_fill_bit~0 .extended_lut = "on";
defparam \A_slow_ld_data_fill_bit~0 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \A_slow_ld_data_fill_bit~0 .shared_arith = "off";

dffeas \A_slow_inst_result[30] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[30]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[30]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[30] .is_wysiwyg = "true";
defparam \A_slow_inst_result[30] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[30]~61 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[30]~q ),
	.dataf(!\A_slow_inst_result[30]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[30]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[30]~61 .extended_lut = "off";
defparam \A_wr_data_unfiltered[30]~61 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[30]~61 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[30]~62 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[30]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[30]~q ),
	.datae(!\A_wr_data_unfiltered[30]~61_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[30]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[30]~62 .extended_lut = "off";
defparam \A_wr_data_unfiltered[30]~62 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[30]~62 .shared_arith = "off";

dffeas \W_wr_data[30] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[30]~62_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[30]~q ),
	.prn(vcc));
defparam \W_wr_data[30] .is_wysiwyg = "true";
defparam \W_wr_data[30] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[30]~14 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[30] ),
	.datab(!\W_wr_data[30]~q ),
	.datac(!\M_alu_result[30]~q ),
	.datad(!\A_wr_data_unfiltered[30]~62_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[30]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[30]~14 .extended_lut = "off";
defparam \D_src1_reg[30]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[30]~14 .shared_arith = "off";

dffeas \E_src1[30] (
	.clk(clk_clk),
	.d(\D_src1_reg[30]~14_combout ),
	.asdata(\E_alu_result[30]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[30]~q ),
	.prn(vcc));
defparam \E_src1[30] .is_wysiwyg = "true";
defparam \E_src1[30] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[1]~10 (
	.dataa(!\E_src1[1]~q ),
	.datab(!\E_src1[0]~q ),
	.datac(!\E_src1[31]~q ),
	.datad(!\E_src1[30]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[1]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[1]~10 .extended_lut = "off";
defparam \E_rot_step1[1]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[1]~10 .shared_arith = "off";

dffeas \M_rot_prestep2[5] (
	.clk(clk_clk),
	.d(\E_rot_step1[1]~10_combout ),
	.asdata(\E_rot_step1[5]~11_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[5]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[5] .is_wysiwyg = "true";
defparam \M_rot_prestep2[5] .power_up = "low";

cyclonev_lcell_comb \M_rot[5]~1 (
	.dataa(!\M_rot_prestep2[13]~q ),
	.datab(!\M_rot_prestep2[5]~q ),
	.datac(!\M_rot_prestep2[29]~q ),
	.datad(!\M_rot_prestep2[21]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~1 .extended_lut = "off";
defparam \M_rot[5]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~1 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_mask[5]~q ),
	.datad(!\M_rot_sel_fill1~q ),
	.datae(!\M_rot[5]~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~1 .extended_lut = "off";
defparam \A_shift_rot_result~1 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~1 .shared_arith = "off";

dffeas \A_shift_rot_result[13] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[13]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[13] .is_wysiwyg = "true";
defparam \A_shift_rot_result[13] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[13]~7 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_mul_result[13]~q ),
	.datac(!\A_shift_rot_result[13]~q ),
	.datad(!\A_ctrl_shift_rot~q ),
	.datae(!\A_wr_data_unfiltered[13]~6_combout ),
	.dataf(!\D_src2_reg[5]~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[13]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[13]~7 .extended_lut = "off";
defparam \D_src2_reg[13]~7 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \D_src2_reg[13]~7 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[13]~92 (
	.dataa(!\M_alu_result[13]~q ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\W_wr_data[13]~q ),
	.datad(!\D_src2_reg[5]~3_combout ),
	.datae(!\D_src2_reg[13]~7_combout ),
	.dataf(!\D_src2_reg[13]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[13]~92_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[13]~92 .extended_lut = "off";
defparam \D_src2_reg[13]~92 .lut_mask = 64'hCF5FFFFFFFFFFFFF;
defparam \D_src2_reg[13]~92 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[13]~0 (
	.dataa(!\E_src2[13]~q ),
	.datab(!\E_src1[13]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[13]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[13]~0 .extended_lut = "off";
defparam \E_logic_result[13]~0 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[13]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ctrl_jmp_indirect_nxt~0 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_iw[11]~q ),
	.datac(!\D_iw[16]~q ),
	.datad(!\Equal171~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_jmp_indirect_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_jmp_indirect_nxt~0 .extended_lut = "off";
defparam \E_ctrl_jmp_indirect_nxt~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \E_ctrl_jmp_indirect_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \E_valid_jmp_indirect~0 (
	.dataa(!\D_valid~combout ),
	.datab(!\E_ctrl_jmp_indirect_nxt~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid_jmp_indirect~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid_jmp_indirect~0 .extended_lut = "off";
defparam \E_valid_jmp_indirect~0 .lut_mask = 64'h7777777777777777;
defparam \E_valid_jmp_indirect~0 .shared_arith = "off";

dffeas E_valid_jmp_indirect(
	.clk(clk_clk),
	.d(\E_valid_jmp_indirect~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_valid_jmp_indirect~q ),
	.prn(vcc));
defparam E_valid_jmp_indirect.is_wysiwyg = "true";
defparam E_valid_jmp_indirect.power_up = "low";

dffeas \D_pc[11] (
	.clk(clk_clk),
	.d(\F_pc[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[11]~q ),
	.prn(vcc));
defparam \D_pc[11] .is_wysiwyg = "true";
defparam \D_pc[11] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[12]~2 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[12] ),
	.datab(!\W_wr_data[12]~q ),
	.datac(!\M_alu_result[12]~q ),
	.datad(!\A_wr_data_unfiltered[12]~9_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[12]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[12]~2 .extended_lut = "off";
defparam \D_src1_reg[12]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[12]~2 .shared_arith = "off";

dffeas \E_src1[12] (
	.clk(clk_clk),
	.d(\D_src1_reg[12]~2_combout ),
	.asdata(\E_alu_result[12]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[12]~q ),
	.prn(vcc));
defparam \E_src1[12] .is_wysiwyg = "true";
defparam \E_src1[12] .power_up = "low";

dffeas \D_pc[10] (
	.clk(clk_clk),
	.d(\F_pc[10]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[10]~q ),
	.prn(vcc));
defparam \D_pc[10] .is_wysiwyg = "true";
defparam \D_pc[10] .power_up = "low";

cyclonev_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~1_sumout ),
	.cout(\Add3~2 ),
	.shareout());
defparam \Add3~1 .extended_lut = "off";
defparam \Add3~1 .lut_mask = 64'h00000000000000FF;
defparam \Add3~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[8] ),
	.datae(gnd),
	.dataf(!\Add3~1_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[0] (
	.clk(clk_clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[0]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[0] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[0] .power_up = "low";

dffeas \D_pc_plus_one[0] (
	.clk(clk_clk),
	.d(\Add3~1_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[0]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[0] .is_wysiwyg = "true";
defparam \D_pc_plus_one[0] .power_up = "low";

cyclonev_lcell_comb \E_ctrl_br_cond_nxt~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_br_cond_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_br_cond_nxt~0 .extended_lut = "off";
defparam \E_ctrl_br_cond_nxt~0 .lut_mask = 64'hAFFF3FFFFFFFFFFF;
defparam \E_ctrl_br_cond_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb D_br_pred_not_taken(
	.dataa(!\D_bht_data[1]~q ),
	.datab(!\E_ctrl_br_cond_nxt~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_br_pred_not_taken~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_br_pred_not_taken.extended_lut = "off";
defparam D_br_pred_not_taken.lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam D_br_pred_not_taken.shared_arith = "off";

dffeas \E_extra_pc[0] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[0]~q ),
	.asdata(\D_pc_plus_one[0]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[0]~q ),
	.prn(vcc));
defparam \E_extra_pc[0] .is_wysiwyg = "true";
defparam \E_extra_pc[0] .power_up = "low";

dffeas E_ctrl_jmp_indirect(
	.clk(clk_clk),
	.d(\E_ctrl_jmp_indirect_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_jmp_indirect~q ),
	.prn(vcc));
defparam E_ctrl_jmp_indirect.is_wysiwyg = "true";
defparam E_ctrl_jmp_indirect.power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[0]~0 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_ctrl_break~q ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_ctrl_jmp_indirect~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[0]~0 .extended_lut = "off";
defparam \M_pipe_flush_waddr[0]~0 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \M_pipe_flush_waddr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[0]~0 (
	.dataa(!\E_src1[2]~q ),
	.datab(!\E_extra_pc[0]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[0]~0 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[0]~0 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[0]~0 .shared_arith = "off";

dffeas \D_pc[0] (
	.clk(clk_clk),
	.d(\F_pc[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[0]~q ),
	.prn(vcc));
defparam \D_pc[0] .is_wysiwyg = "true";
defparam \D_pc[0] .power_up = "low";

dffeas \E_pc[0] (
	.clk(clk_clk),
	.d(\D_pc[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[0]~q ),
	.prn(vcc));
defparam \E_pc[0] .is_wysiwyg = "true";
defparam \E_pc[0] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[0]~1 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_ctrl_jmp_indirect~q ),
	.datac(!\E_ctrl_crst~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[0]~1 .extended_lut = "off";
defparam \M_pipe_flush_waddr[0]~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \M_pipe_flush_waddr[0]~1 .shared_arith = "off";

dffeas \M_pipe_flush_waddr[0] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[0]~0_combout ),
	.asdata(\E_pc[0]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[0]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[0] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[0] .power_up = "low";

dffeas D_kill(
	.clk(clk_clk),
	.d(\F_kill~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_kill~q ),
	.prn(vcc));
defparam D_kill.is_wysiwyg = "true";
defparam D_kill.power_up = "low";

cyclonev_lcell_comb \F_ctrl_br~0 (
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[1]~3_combout ),
	.datac(!\F_iw[2]~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_br~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_br~0 .extended_lut = "off";
defparam \F_ctrl_br~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \F_ctrl_br~0 .shared_arith = "off";

dffeas D_ctrl_br(
	.clk(clk_clk),
	.d(\F_ctrl_br~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_br~q ),
	.prn(vcc));
defparam D_ctrl_br.is_wysiwyg = "true";
defparam D_ctrl_br.power_up = "low";

cyclonev_lcell_comb \F_ctrl_br_uncond~0 (
	.dataa(!\F_iw[0]~9_combout ),
	.datab(!\F_iw[5]~1_combout ),
	.datac(!\F_iw[3]~2_combout ),
	.datad(!\F_iw[1]~3_combout ),
	.datae(!\F_iw[4]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ctrl_br_uncond~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ctrl_br_uncond~0 .extended_lut = "off";
defparam \F_ctrl_br_uncond~0 .lut_mask = 64'hFFFFFEFFFFFFFEFF;
defparam \F_ctrl_br_uncond~0 .shared_arith = "off";

dffeas D_ctrl_br_uncond(
	.clk(clk_clk),
	.d(\F_ctrl_br_uncond~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ctrl_br_uncond~q ),
	.prn(vcc));
defparam D_ctrl_br_uncond.is_wysiwyg = "true";
defparam D_ctrl_br_uncond.power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[2]~1 (
	.dataa(!\D_issue~q ),
	.datab(!\D_bht_data[1]~q ),
	.datac(!\D_iw_valid~q ),
	.datad(!\D_kill~q ),
	.datae(!\D_ctrl_br~q ),
	.dataf(!\D_ctrl_br_uncond~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[2]~1 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[2]~1 .lut_mask = 64'hFFFDFFFFFFFFFFFF;
defparam \F_ic_data_rd_addr_nxt[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[0]~2 (
	.dataa(!\D_pc[0]~q ),
	.datab(!\D_br_taken_waddr_partial[0]~q ),
	.datac(!\Add3~1_sumout ),
	.datad(!\D_iw[6]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[0]~2 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[0]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[0]~3 (
	.dataa(!\E_src1[2]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[0]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[0]~3 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[0]~3 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_data_rd_addr_nxt[0]~3 .shared_arith = "off";

dffeas \F_pc[0] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[0]~q ),
	.prn(vcc));
defparam \F_pc[0] .is_wysiwyg = "true";
defparam \F_pc[0] .power_up = "low";

cyclonev_lcell_comb \Add3~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~45_sumout ),
	.cout(\Add3~46 ),
	.shareout());
defparam \Add3~45 .extended_lut = "off";
defparam \Add3~45 .lut_mask = 64'h00000000000000FF;
defparam \Add3~45 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[9] ),
	.datae(gnd),
	.dataf(!\Add3~45_sumout ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[1] (
	.clk(clk_clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[1]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[1] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[1] .power_up = "low";

dffeas \D_pc_plus_one[1] (
	.clk(clk_clk),
	.d(\Add3~45_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[1]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[1] .is_wysiwyg = "true";
defparam \D_pc_plus_one[1] .power_up = "low";

dffeas \E_extra_pc[1] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[1]~q ),
	.asdata(\D_pc_plus_one[1]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[1]~q ),
	.prn(vcc));
defparam \E_extra_pc[1] .is_wysiwyg = "true";
defparam \E_extra_pc[1] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[1]~1 (
	.dataa(!\E_src1[3]~q ),
	.datab(!\E_extra_pc[1]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[1]~1 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[1]~1 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[1]~1 .shared_arith = "off";

dffeas \D_pc[1] (
	.clk(clk_clk),
	.d(\F_pc[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[1]~q ),
	.prn(vcc));
defparam \D_pc[1] .is_wysiwyg = "true";
defparam \D_pc[1] .power_up = "low";

dffeas \E_pc[1] (
	.clk(clk_clk),
	.d(\D_pc[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[1]~q ),
	.prn(vcc));
defparam \E_pc[1] .is_wysiwyg = "true";
defparam \E_pc[1] .power_up = "low";

dffeas \M_pipe_flush_waddr[1] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[1]~1_combout ),
	.asdata(\E_pc[1]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[1]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[1] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[1] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[1]~4 (
	.dataa(!\D_pc[1]~q ),
	.datab(!\D_br_taken_waddr_partial[1]~q ),
	.datac(!\Add3~45_sumout ),
	.datad(!\D_iw[7]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[1]~4 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[1]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[1]~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[1]~5 (
	.dataa(!\E_src1[3]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[1]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[1]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[1]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[1]~5 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[1]~5 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_data_rd_addr_nxt[1]~5 .shared_arith = "off";

dffeas \F_pc[1] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[1]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[1]~q ),
	.prn(vcc));
defparam \F_pc[1] .is_wysiwyg = "true";
defparam \F_pc[1] .power_up = "low";

cyclonev_lcell_comb \Add3~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~41_sumout ),
	.cout(\Add3~42 ),
	.shareout());
defparam \Add3~41 .extended_lut = "off";
defparam \Add3~41 .lut_mask = 64'h00000000000000FF;
defparam \Add3~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[10] ),
	.datae(gnd),
	.dataf(!\Add3~41_sumout ),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[2] (
	.clk(clk_clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[2]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[2] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[2] .power_up = "low";

dffeas \D_pc_plus_one[2] (
	.clk(clk_clk),
	.d(\Add3~41_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[2]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[2] .is_wysiwyg = "true";
defparam \D_pc_plus_one[2] .power_up = "low";

dffeas \E_extra_pc[2] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[2]~q ),
	.asdata(\D_pc_plus_one[2]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[2]~q ),
	.prn(vcc));
defparam \E_extra_pc[2] .is_wysiwyg = "true";
defparam \E_extra_pc[2] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[2]~2 (
	.dataa(!\E_src1[4]~q ),
	.datab(!\E_extra_pc[2]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[2]~2 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[2]~2 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[2]~2 .shared_arith = "off";

dffeas \D_pc[2] (
	.clk(clk_clk),
	.d(\F_pc[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[2]~q ),
	.prn(vcc));
defparam \D_pc[2] .is_wysiwyg = "true";
defparam \D_pc[2] .power_up = "low";

dffeas \E_pc[2] (
	.clk(clk_clk),
	.d(\D_pc[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[2]~q ),
	.prn(vcc));
defparam \E_pc[2] .is_wysiwyg = "true";
defparam \E_pc[2] .power_up = "low";

dffeas \M_pipe_flush_waddr[2] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[2]~2_combout ),
	.asdata(\E_pc[2]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[2]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[2] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[2] .power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[2]~6 (
	.dataa(!\D_pc[2]~q ),
	.datab(!\D_br_taken_waddr_partial[2]~q ),
	.datac(!\Add3~41_sumout ),
	.datad(!\D_iw[8]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[2]~6 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[2]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_data_rd_addr_nxt[2]~6 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[2]~7 (
	.dataa(!\E_src1[4]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[2]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[2]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[2]~7 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[2]~7 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_data_rd_addr_nxt[2]~7 .shared_arith = "off";

dffeas \F_pc[2] (
	.clk(clk_clk),
	.d(\F_ic_data_rd_addr_nxt[2]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[2]~q ),
	.prn(vcc));
defparam \F_pc[2] .is_wysiwyg = "true";
defparam \F_pc[2] .power_up = "low";

cyclonev_lcell_comb \Add3~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~37_sumout ),
	.cout(\Add3~38 ),
	.shareout());
defparam \Add3~37 .extended_lut = "off";
defparam \Add3~37 .lut_mask = 64'h00000000000000FF;
defparam \Add3~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[11] ),
	.datae(gnd),
	.dataf(!\Add3~37_sumout ),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[3] (
	.clk(clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[3]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[3] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[3] .power_up = "low";

dffeas \D_pc_plus_one[3] (
	.clk(clk_clk),
	.d(\Add3~37_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[3]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[3] .is_wysiwyg = "true";
defparam \D_pc_plus_one[3] .power_up = "low";

dffeas \E_extra_pc[3] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[3]~q ),
	.asdata(\D_pc_plus_one[3]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[3]~q ),
	.prn(vcc));
defparam \E_extra_pc[3] .is_wysiwyg = "true";
defparam \E_extra_pc[3] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[3]~3 (
	.dataa(!\E_src1[5]~q ),
	.datab(!\E_extra_pc[3]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[3]~3 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[3]~3 .lut_mask = 64'h53FF53FF53FF53FF;
defparam \M_pipe_flush_waddr_nxt[3]~3 .shared_arith = "off";

dffeas \D_pc[3] (
	.clk(clk_clk),
	.d(\F_pc[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[3]~q ),
	.prn(vcc));
defparam \D_pc[3] .is_wysiwyg = "true";
defparam \D_pc[3] .power_up = "low";

dffeas \E_pc[3] (
	.clk(clk_clk),
	.d(\D_pc[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[3]~q ),
	.prn(vcc));
defparam \E_pc[3] .is_wysiwyg = "true";
defparam \E_pc[3] .power_up = "low";

dffeas \M_pipe_flush_waddr[3] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[3]~3_combout ),
	.asdata(\E_pc[3]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[3]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[3] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[3] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[0]~0 (
	.dataa(!\D_pc[3]~q ),
	.datab(!\D_br_taken_waddr_partial[3]~q ),
	.datac(!\Add3~37_sumout ),
	.datad(!\D_iw[9]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[0]~0 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[0]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[0]~1 (
	.dataa(!\E_src1[5]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[3]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[0]~1 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[0]~1 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[0]~1 .shared_arith = "off";

dffeas \F_pc[3] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[3]~q ),
	.prn(vcc));
defparam \F_pc[3] .is_wysiwyg = "true";
defparam \F_pc[3] .power_up = "low";

cyclonev_lcell_comb \Add3~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~33_sumout ),
	.cout(\Add3~34 ),
	.shareout());
defparam \Add3~33 .extended_lut = "off";
defparam \Add3~33 .lut_mask = 64'h00000000000000FF;
defparam \Add3~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[12] ),
	.datae(gnd),
	.dataf(!\Add3~33_sumout ),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[4] (
	.clk(clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[4]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[4] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[4] .power_up = "low";

dffeas \D_pc_plus_one[4] (
	.clk(clk_clk),
	.d(\Add3~33_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[4]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[4] .is_wysiwyg = "true";
defparam \D_pc_plus_one[4] .power_up = "low";

dffeas \E_extra_pc[4] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[4]~q ),
	.asdata(\D_pc_plus_one[4]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[4]~q ),
	.prn(vcc));
defparam \E_extra_pc[4] .is_wysiwyg = "true";
defparam \E_extra_pc[4] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[4]~4 (
	.dataa(!\E_src1[6]~q ),
	.datab(!\E_extra_pc[4]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[4]~4 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[4]~4 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[4]~4 .shared_arith = "off";

dffeas \D_pc[4] (
	.clk(clk_clk),
	.d(\F_pc[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[4]~q ),
	.prn(vcc));
defparam \D_pc[4] .is_wysiwyg = "true";
defparam \D_pc[4] .power_up = "low";

dffeas \E_pc[4] (
	.clk(clk_clk),
	.d(\D_pc[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[4]~q ),
	.prn(vcc));
defparam \E_pc[4] .is_wysiwyg = "true";
defparam \E_pc[4] .power_up = "low";

dffeas \M_pipe_flush_waddr[4] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[4]~4_combout ),
	.asdata(\E_pc[4]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[4]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[4] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[4] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[1]~2 (
	.dataa(!\D_pc[4]~q ),
	.datab(!\D_br_taken_waddr_partial[4]~q ),
	.datac(!\Add3~33_sumout ),
	.datad(!\D_iw[10]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[1]~2 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[1]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[1]~3 (
	.dataa(!\E_src1[6]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[4]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[1]~3 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[1]~3 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[1]~3 .shared_arith = "off";

dffeas \F_pc[4] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[1]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[4]~q ),
	.prn(vcc));
defparam \F_pc[4] .is_wysiwyg = "true";
defparam \F_pc[4] .power_up = "low";

cyclonev_lcell_comb \Add3~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~29_sumout ),
	.cout(\Add3~30 ),
	.shareout());
defparam \Add3~29 .extended_lut = "off";
defparam \Add3~29 .lut_mask = 64'h00000000000000FF;
defparam \Add3~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[13] ),
	.datae(gnd),
	.dataf(!\Add3~29_sumout ),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[5] (
	.clk(clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[5]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[5] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[5] .power_up = "low";

dffeas \D_pc_plus_one[5] (
	.clk(clk_clk),
	.d(\Add3~29_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[5]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[5] .is_wysiwyg = "true";
defparam \D_pc_plus_one[5] .power_up = "low";

dffeas \E_extra_pc[5] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[5]~q ),
	.asdata(\D_pc_plus_one[5]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[5]~q ),
	.prn(vcc));
defparam \E_extra_pc[5] .is_wysiwyg = "true";
defparam \E_extra_pc[5] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[5]~5 (
	.dataa(!\E_src1[7]~q ),
	.datab(!\E_extra_pc[5]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[5]~5 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[5]~5 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[5]~5 .shared_arith = "off";

dffeas \D_pc[5] (
	.clk(clk_clk),
	.d(\F_pc[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[5]~q ),
	.prn(vcc));
defparam \D_pc[5] .is_wysiwyg = "true";
defparam \D_pc[5] .power_up = "low";

dffeas \E_pc[5] (
	.clk(clk_clk),
	.d(\D_pc[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[5]~q ),
	.prn(vcc));
defparam \E_pc[5] .is_wysiwyg = "true";
defparam \E_pc[5] .power_up = "low";

dffeas \M_pipe_flush_waddr[5] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[5]~5_combout ),
	.asdata(\E_pc[5]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[5]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[5] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[5] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[2]~4 (
	.dataa(!\D_pc[5]~q ),
	.datab(!\D_br_taken_waddr_partial[5]~q ),
	.datac(!\Add3~29_sumout ),
	.datad(!\D_iw[11]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[2]~4 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[2]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[2]~5 (
	.dataa(!\E_src1[7]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[5]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[2]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[2]~5 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[2]~5 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[2]~5 .shared_arith = "off";

dffeas \F_pc[5] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[2]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[5]~q ),
	.prn(vcc));
defparam \F_pc[5] .is_wysiwyg = "true";
defparam \F_pc[5] .power_up = "low";

cyclonev_lcell_comb \Add3~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~25_sumout ),
	.cout(\Add3~26 ),
	.shareout());
defparam \Add3~25 .extended_lut = "off";
defparam \Add3~25 .lut_mask = 64'h00000000000000FF;
defparam \Add3~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[14] ),
	.datae(gnd),
	.dataf(!\Add3~25_sumout ),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[6] (
	.clk(clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[6]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[6] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[6] .power_up = "low";

dffeas \D_pc_plus_one[6] (
	.clk(clk_clk),
	.d(\Add3~25_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[6]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[6] .is_wysiwyg = "true";
defparam \D_pc_plus_one[6] .power_up = "low";

dffeas \E_extra_pc[6] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[6]~q ),
	.asdata(\D_pc_plus_one[6]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[6]~q ),
	.prn(vcc));
defparam \E_extra_pc[6] .is_wysiwyg = "true";
defparam \E_extra_pc[6] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[6]~6 (
	.dataa(!\E_src1[8]~q ),
	.datab(!\E_extra_pc[6]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[6]~6 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[6]~6 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[6]~6 .shared_arith = "off";

dffeas \D_pc[6] (
	.clk(clk_clk),
	.d(\F_pc[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[6]~q ),
	.prn(vcc));
defparam \D_pc[6] .is_wysiwyg = "true";
defparam \D_pc[6] .power_up = "low";

dffeas \E_pc[6] (
	.clk(clk_clk),
	.d(\D_pc[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[6]~q ),
	.prn(vcc));
defparam \E_pc[6] .is_wysiwyg = "true";
defparam \E_pc[6] .power_up = "low";

dffeas \M_pipe_flush_waddr[6] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[6]~6_combout ),
	.asdata(\E_pc[6]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[6]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[6] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[6] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~6 (
	.dataa(!\D_pc[6]~q ),
	.datab(!\D_br_taken_waddr_partial[6]~q ),
	.datac(!\Add3~25_sumout ),
	.datad(!\D_iw[12]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~6 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[3]~6 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[3]~7 (
	.dataa(!\E_src1[8]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[6]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[3]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[3]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[3]~7 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[3]~7 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[3]~7 .shared_arith = "off";

dffeas \F_pc[6] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[3]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[6]~q ),
	.prn(vcc));
defparam \F_pc[6] .is_wysiwyg = "true";
defparam \F_pc[6] .power_up = "low";

cyclonev_lcell_comb \Add3~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~21_sumout ),
	.cout(\Add3~22 ),
	.shareout());
defparam \Add3~21 .extended_lut = "off";
defparam \Add3~21 .lut_mask = 64'h00000000000000FF;
defparam \Add3~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[15] ),
	.datae(gnd),
	.dataf(!\Add3~21_sumout ),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[7] (
	.clk(clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[7]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[7] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[7] .power_up = "low";

dffeas \D_pc_plus_one[7] (
	.clk(clk_clk),
	.d(\Add3~21_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[7]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[7] .is_wysiwyg = "true";
defparam \D_pc_plus_one[7] .power_up = "low";

dffeas \E_extra_pc[7] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[7]~q ),
	.asdata(\D_pc_plus_one[7]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[7]~q ),
	.prn(vcc));
defparam \E_extra_pc[7] .is_wysiwyg = "true";
defparam \E_extra_pc[7] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[7]~7 (
	.dataa(!\E_src1[9]~q ),
	.datab(!\E_extra_pc[7]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[7]~7 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[7]~7 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[7]~7 .shared_arith = "off";

dffeas \D_pc[7] (
	.clk(clk_clk),
	.d(\F_pc[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[7]~q ),
	.prn(vcc));
defparam \D_pc[7] .is_wysiwyg = "true";
defparam \D_pc[7] .power_up = "low";

dffeas \E_pc[7] (
	.clk(clk_clk),
	.d(\D_pc[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[7]~q ),
	.prn(vcc));
defparam \E_pc[7] .is_wysiwyg = "true";
defparam \E_pc[7] .power_up = "low";

dffeas \M_pipe_flush_waddr[7] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[7]~7_combout ),
	.asdata(\E_pc[7]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[7]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[7] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[7] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[4]~8 (
	.dataa(!\D_pc[7]~q ),
	.datab(!\D_br_taken_waddr_partial[7]~q ),
	.datac(!\Add3~21_sumout ),
	.datad(!\D_iw[13]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[4]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[4]~8 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[4]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[4]~8 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[4]~9 (
	.dataa(!\E_src1[9]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[7]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[4]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[4]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[4]~9 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[4]~9 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[4]~9 .shared_arith = "off";

dffeas \F_pc[7] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[4]~9_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[7]~q ),
	.prn(vcc));
defparam \F_pc[7] .is_wysiwyg = "true";
defparam \F_pc[7] .power_up = "low";

cyclonev_lcell_comb \Add3~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~17_sumout ),
	.cout(\Add3~18 ),
	.shareout());
defparam \Add3~17 .extended_lut = "off";
defparam \Add3~17 .lut_mask = 64'h00000000000000FF;
defparam \Add3~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[16] ),
	.datae(gnd),
	.dataf(!\Add3~17_sumout ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[8] (
	.clk(clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[8]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[8] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[8] .power_up = "low";

dffeas \D_pc_plus_one[8] (
	.clk(clk_clk),
	.d(\Add3~17_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[8]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[8] .is_wysiwyg = "true";
defparam \D_pc_plus_one[8] .power_up = "low";

dffeas \E_extra_pc[8] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[8]~q ),
	.asdata(\D_pc_plus_one[8]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[8]~q ),
	.prn(vcc));
defparam \E_extra_pc[8] .is_wysiwyg = "true";
defparam \E_extra_pc[8] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[8]~8 (
	.dataa(!\E_src1[10]~q ),
	.datab(!\E_extra_pc[8]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[0]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[8]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[8]~8 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[8]~8 .lut_mask = 64'hF737F737F737F737;
defparam \M_pipe_flush_waddr_nxt[8]~8 .shared_arith = "off";

dffeas \D_pc[8] (
	.clk(clk_clk),
	.d(\F_pc[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[8]~q ),
	.prn(vcc));
defparam \D_pc[8] .is_wysiwyg = "true";
defparam \D_pc[8] .power_up = "low";

dffeas \E_pc[8] (
	.clk(clk_clk),
	.d(\D_pc[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[8]~q ),
	.prn(vcc));
defparam \E_pc[8] .is_wysiwyg = "true";
defparam \E_pc[8] .power_up = "low";

dffeas \M_pipe_flush_waddr[8] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[8]~8_combout ),
	.asdata(\E_pc[8]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[8]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[8] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[8] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[5]~10 (
	.dataa(!\D_pc[8]~q ),
	.datab(!\D_br_taken_waddr_partial[8]~q ),
	.datac(!\Add3~17_sumout ),
	.datad(!\D_iw[14]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[5]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[5]~10 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[5]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[5]~10 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[5]~11 (
	.dataa(!\E_src1[10]~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[8]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[5]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[5]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[5]~11 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[5]~11 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[5]~11 .shared_arith = "off";

dffeas \F_pc[8] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[5]~11_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[8]~q ),
	.prn(vcc));
defparam \F_pc[8] .is_wysiwyg = "true";
defparam \F_pc[8] .power_up = "low";

cyclonev_lcell_comb \Add3~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~13_sumout ),
	.cout(\Add3~14 ),
	.shareout());
defparam \Add3~13 .extended_lut = "off";
defparam \Add3~13 .lut_mask = 64'h00000000000000FF;
defparam \Add3~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[17] ),
	.datae(gnd),
	.dataf(!\Add3~13_sumout ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[9] (
	.clk(clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[9]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[9] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[9] .power_up = "low";

dffeas \D_pc_plus_one[9] (
	.clk(clk_clk),
	.d(\Add3~13_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[9]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[9] .is_wysiwyg = "true";
defparam \D_pc_plus_one[9] .power_up = "low";

dffeas \E_extra_pc[9] (
	.clk(clk_clk),
	.d(\D_br_taken_waddr_partial[9]~q ),
	.asdata(\D_pc_plus_one[9]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[9]~q ),
	.prn(vcc));
defparam \E_extra_pc[9] .is_wysiwyg = "true";
defparam \E_extra_pc[9] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[9]~9 (
	.dataa(!\E_src1[11]~q ),
	.datab(!\E_extra_pc[9]~q ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_ctrl_jmp_indirect~q ),
	.datae(!\M_pipe_flush_waddr[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[9]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[9]~9 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[9]~9 .lut_mask = 64'hF7FFFFF7F7FFFFF7;
defparam \M_pipe_flush_waddr_nxt[9]~9 .shared_arith = "off";

dffeas \D_pc[9] (
	.clk(clk_clk),
	.d(\F_pc[9]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc[9]~q ),
	.prn(vcc));
defparam \D_pc[9] .is_wysiwyg = "true";
defparam \D_pc[9] .power_up = "low";

dffeas \E_pc[9] (
	.clk(clk_clk),
	.d(\D_pc[9]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[9]~q ),
	.prn(vcc));
defparam \E_pc[9] .is_wysiwyg = "true";
defparam \E_pc[9] .power_up = "low";

dffeas \M_pipe_flush_waddr[9] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[9]~9_combout ),
	.asdata(\E_pc[9]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[9]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[9] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[9] .power_up = "low";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[6]~12 (
	.dataa(!\D_pc[9]~q ),
	.datab(!\D_br_taken_waddr_partial[9]~q ),
	.datac(!\Add3~13_sumout ),
	.datad(!\D_iw[15]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[6]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[6]~12 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[6]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_ic_tag_rd_addr_nxt[6]~12 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_tag_rd_addr_nxt[6]~13 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\E_src1[11]~q ),
	.datac(!\E_valid_jmp_indirect~q ),
	.datad(!\M_pipe_flush_waddr[9]~q ),
	.datae(!\F_ic_tag_rd_addr_nxt[6]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_tag_rd_addr_nxt[6]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_tag_rd_addr_nxt[6]~13 .extended_lut = "off";
defparam \F_ic_tag_rd_addr_nxt[6]~13 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \F_ic_tag_rd_addr_nxt[6]~13 .shared_arith = "off";

dffeas \F_pc[9] (
	.clk(clk_clk),
	.d(\F_ic_tag_rd_addr_nxt[6]~13_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\F_pc[9]~q ),
	.prn(vcc));
defparam \F_pc[9] .is_wysiwyg = "true";
defparam \F_pc[9] .power_up = "low";

cyclonev_lcell_comb \Add3~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~9_sumout ),
	.cout(\Add3~10 ),
	.shareout());
defparam \Add3~9 .extended_lut = "off";
defparam \Add3~9 .lut_mask = 64'h00000000000000FF;
defparam \Add3~9 .shared_arith = "off";

dffeas \D_pc_plus_one[10] (
	.clk(clk_clk),
	.d(\Add3~9_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[10]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[10] .is_wysiwyg = "true";
defparam \D_pc_plus_one[10] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000000000000000;
defparam \Add0~5 .shared_arith = "off";

dffeas \D_br_taken_waddr_partial[10] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_br_taken_waddr_partial[10]~q ),
	.prn(vcc));
defparam \D_br_taken_waddr_partial[10] .is_wysiwyg = "true";
defparam \D_br_taken_waddr_partial[10] .power_up = "low";

cyclonev_lcell_comb \Add1~1 (
	.dataa(!\D_iw[18]~q ),
	.datab(!\D_pc_plus_one[10]~q ),
	.datac(!\D_br_taken_waddr_partial[10]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h9696969696969696;
defparam \Add1~1 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~0 (
	.dataa(!\D_pc[10]~q ),
	.datab(!\Add1~1_combout ),
	.datac(!\Add3~9_sumout ),
	.datad(!\D_iw[16]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~0 .extended_lut = "off";
defparam \F_pc_nxt~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~1 (
	.dataa(!\E_src1[12]~q ),
	.datab(!\E_valid_jmp_indirect~q ),
	.datac(!\F_pc_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~1 .extended_lut = "off";
defparam \F_pc_nxt~1 .lut_mask = 64'h4747474747474747;
defparam \F_pc_nxt~1 .shared_arith = "off";

dffeas \E_pc[10] (
	.clk(clk_clk),
	.d(\D_pc[10]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[10]~q ),
	.prn(vcc));
defparam \E_pc[10] .is_wysiwyg = "true";
defparam \E_pc[10] .power_up = "low";

dffeas \E_extra_pc[10] (
	.clk(clk_clk),
	.d(\Add1~1_combout ),
	.asdata(\D_pc_plus_one[10]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[10]~q ),
	.prn(vcc));
defparam \E_extra_pc[10] .is_wysiwyg = "true";
defparam \E_extra_pc[10] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[10]~10 (
	.dataa(!\E_extra_pc[10]~q ),
	.datab(!\E_ctrl_break~q ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_ctrl_crst~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[10]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[10]~10 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[10]~10 .lut_mask = 64'hFFFBFFFBFFFBFFFB;
defparam \M_pipe_flush_waddr_nxt[10]~10 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[10]~11 (
	.dataa(!\E_hbreak_req~combout ),
	.datab(!\E_src1[12]~q ),
	.datac(!\E_ctrl_jmp_indirect~q ),
	.datad(!\E_pc[10]~q ),
	.datae(!\M_pipe_flush_waddr_nxt[10]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[10]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[10]~11 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[10]~11 .lut_mask = 64'hFFDEFFFFFFDEFFFF;
defparam \M_pipe_flush_waddr_nxt[10]~11 .shared_arith = "off";

dffeas \M_pipe_flush_waddr[10] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[10]~11_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[10]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[10] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[10] .power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_waddr[10]~_wirecell (
	.dataa(!\M_pipe_flush_waddr[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr[10]~_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr[10]~_wirecell .extended_lut = "off";
defparam \M_pipe_flush_waddr[10]~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \M_pipe_flush_waddr[10]~_wirecell .shared_arith = "off";

dffeas \F_pc[10] (
	.clk(clk_clk),
	.d(\F_pc_nxt~1_combout ),
	.asdata(\M_pipe_flush_waddr[10]~_wirecell_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\M_pipe_flush~q ),
	.ena(!\F_stall~combout ),
	.q(\F_pc[10]~q ),
	.prn(vcc));
defparam \F_pc[10] .is_wysiwyg = "true";
defparam \F_pc[10] .power_up = "low";

cyclonev_lcell_comb \F_ic_valid~4 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[3] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[5] ),
	.datac(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[4] ),
	.datad(!\F_pc[0]~q ),
	.datae(!\F_pc[1]~q ),
	.dataf(!\F_pc[2]~q ),
	.datag(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[2] ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_valid~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_valid~4 .extended_lut = "on";
defparam \F_ic_valid~4 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \F_ic_valid~4 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_valid~0 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[7] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[9] ),
	.datac(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[8] ),
	.datad(!\F_pc[2]~q ),
	.datae(!\F_pc[1]~q ),
	.dataf(!\F_ic_valid~4_combout ),
	.datag(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[6] ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_valid~0 .extended_lut = "on";
defparam \F_ic_valid~0 .lut_mask = 64'hFAFCFAFCFAFCFAFC;
defparam \F_ic_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_hit~0 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[0] ),
	.datab(!\F_pc[10]~q ),
	.datac(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[1] ),
	.datad(!\F_pc[11]~q ),
	.datae(!\F_ic_valid~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_hit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_hit~0 .extended_lut = "off";
defparam \F_ic_hit~0 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \F_ic_hit~0 .shared_arith = "off";

dffeas D_iw_valid(
	.clk(clk_clk),
	.d(\F_ic_hit~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw_valid~q ),
	.prn(vcc));
defparam D_iw_valid.is_wysiwyg = "true";
defparam D_iw_valid.power_up = "low";

cyclonev_lcell_comb \D_br_pred_taken~0 (
	.dataa(!\D_bht_data[1]~q ),
	.datab(!\D_ctrl_br~q ),
	.datac(!\D_ctrl_br_uncond~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_br_pred_taken~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_br_pred_taken~0 .extended_lut = "off";
defparam \D_br_pred_taken~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \D_br_pred_taken~0 .shared_arith = "off";

cyclonev_lcell_comb \F_kill~2 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\Equal171~0_combout ),
	.datac(!\D_iw[16]~q ),
	.datad(!\D_iw[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_kill~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_kill~2 .extended_lut = "off";
defparam \F_kill~2 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \F_kill~2 .shared_arith = "off";

cyclonev_lcell_comb \F_kill~0 (
	.dataa(!\D_iw[1]~q ),
	.datab(!\D_issue~q ),
	.datac(!\Equal105~0_combout ),
	.datad(!\D_br_pred_taken~0_combout ),
	.datae(!\F_kill~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_kill~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_kill~0 .extended_lut = "off";
defparam \F_kill~0 .lut_mask = 64'hBFFFFFFFBFFFFFFF;
defparam \F_kill~0 .shared_arith = "off";

cyclonev_lcell_comb \F_kill~1 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_iw_valid~q ),
	.datac(!\D_kill~q ),
	.datad(!\E_valid_jmp_indirect~q ),
	.datae(!\F_kill~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_kill~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_kill~1 .extended_lut = "off";
defparam \F_kill~1 .lut_mask = 64'hFEFFFFFFFEFFFFFF;
defparam \F_kill~1 .shared_arith = "off";

cyclonev_lcell_comb F_issue(
	.dataa(!\F_kill~1_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[0] ),
	.datac(!\F_pc[10]~q ),
	.datad(!\embedded_system_nios2_qsys_0_ic_tag|the_altsyncram|auto_generated|q_b[1] ),
	.datae(!\F_pc[11]~q ),
	.dataf(!\F_ic_valid~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_issue~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_issue.extended_lut = "off";
defparam F_issue.lut_mask = 64'hBEEBEBBEFFFFFFFF;
defparam F_issue.shared_arith = "off";

dffeas D_issue(
	.clk(clk_clk),
	.d(\F_issue~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_issue~q ),
	.prn(vcc));
defparam D_issue.is_wysiwyg = "true";
defparam D_issue.power_up = "low";

cyclonev_lcell_comb \F_ic_data_rd_addr_nxt[2]~0 (
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\D_issue~q ),
	.datac(!\D_iw_valid~q ),
	.datad(!\D_kill~q ),
	.datae(!\D_br_pred_taken~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_data_rd_addr_nxt[2]~0 .extended_lut = "off";
defparam \F_ic_data_rd_addr_nxt[2]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \F_ic_data_rd_addr_nxt[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~2 (
	.dataa(!\D_pc[11]~q ),
	.datab(!\Add1~0_combout ),
	.datac(!\Add3~5_sumout ),
	.datad(!\D_iw[17]~q ),
	.datae(!\F_ic_data_rd_addr_nxt[2]~0_combout ),
	.dataf(!\F_ic_data_rd_addr_nxt[2]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~2 .extended_lut = "off";
defparam \F_pc_nxt~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \F_pc_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \F_pc_nxt~3 (
	.dataa(!\E_src1[13]~q ),
	.datab(!\E_valid_jmp_indirect~q ),
	.datac(!\F_pc_nxt~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_pc_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_pc_nxt~3 .extended_lut = "off";
defparam \F_pc_nxt~3 .lut_mask = 64'h4747474747474747;
defparam \F_pc_nxt~3 .shared_arith = "off";

cyclonev_lcell_comb \M_pipe_flush_waddr_nxt[11]~12 (
	.dataa(!\E_src1[13]~q ),
	.datab(!\E_extra_pc[11]~q ),
	.datac(!\E_ctrl_exception~q ),
	.datad(!\E_ctrl_jmp_indirect~q ),
	.datae(!\M_pipe_flush_waddr[0]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_waddr_nxt[11]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_waddr_nxt[11]~12 .extended_lut = "off";
defparam \M_pipe_flush_waddr_nxt[11]~12 .lut_mask = 64'hF7FFFFF7F7FFFFF7;
defparam \M_pipe_flush_waddr_nxt[11]~12 .shared_arith = "off";

dffeas \E_pc[11] (
	.clk(clk_clk),
	.d(\D_pc[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_pc[11]~q ),
	.prn(vcc));
defparam \E_pc[11] .is_wysiwyg = "true";
defparam \E_pc[11] .power_up = "low";

dffeas \M_pipe_flush_waddr[11] (
	.clk(clk_clk),
	.d(\M_pipe_flush_waddr_nxt[11]~12_combout ),
	.asdata(\E_pc[11]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_pipe_flush_waddr[0]~1_combout ),
	.sload(\E_hbreak_req~combout ),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush_waddr[11]~q ),
	.prn(vcc));
defparam \M_pipe_flush_waddr[11] .is_wysiwyg = "true";
defparam \M_pipe_flush_waddr[11] .power_up = "low";

dffeas \F_pc[11] (
	.clk(clk_clk),
	.d(\F_pc_nxt~3_combout ),
	.asdata(\M_pipe_flush_waddr[11]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\M_pipe_flush~q ),
	.ena(!\F_stall~combout ),
	.q(\F_pc[11]~q ),
	.prn(vcc));
defparam \F_pc[11] .is_wysiwyg = "true";
defparam \F_pc[11] .power_up = "low";

cyclonev_lcell_comb \Add3~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\F_pc[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add3~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add3~5_sumout ),
	.cout(),
	.shareout());
defparam \Add3~5 .extended_lut = "off";
defparam \Add3~5 .lut_mask = 64'h00000000000000FF;
defparam \Add3~5 .shared_arith = "off";

dffeas \D_pc_plus_one[11] (
	.clk(clk_clk),
	.d(\Add3~5_sumout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_pc_plus_one[11]~q ),
	.prn(vcc));
defparam \D_pc_plus_one[11] .is_wysiwyg = "true";
defparam \D_pc_plus_one[11] .power_up = "low";

cyclonev_lcell_comb \Add1~0 (
	.dataa(!\D_iw[19]~q ),
	.datab(!\D_pc_plus_one[11]~q ),
	.datac(!\D_iw[18]~q ),
	.datad(!\D_pc_plus_one[10]~q ),
	.datae(!\D_br_taken_waddr_partial[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add1~0 .extended_lut = "off";
defparam \Add1~0 .lut_mask = 64'h9669699696696996;
defparam \Add1~0 .shared_arith = "off";

dffeas \E_extra_pc[11] (
	.clk(clk_clk),
	.d(\Add1~0_combout ),
	.asdata(\D_pc_plus_one[11]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\D_br_pred_not_taken~combout ),
	.ena(\A_stall~combout ),
	.q(\E_extra_pc[11]~q ),
	.prn(vcc));
defparam \E_extra_pc[11] .is_wysiwyg = "true";
defparam \E_extra_pc[11] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[13]~2 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[13]~0_combout ),
	.datac(!\E_ctrl_retaddr~q ),
	.datad(!\E_extra_pc[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[13]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[13]~2 .extended_lut = "off";
defparam \E_alu_result[13]~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[13]~2 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[13]~128 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[13] ),
	.datad(!\D_src2_reg[13]~92_combout ),
	.datae(!\D_src2_reg[5]~2_combout ),
	.dataf(!\E_alu_result[13]~2_combout ),
	.datag(!\Add17~41_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[13]~128_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[13]~128 .extended_lut = "on";
defparam \D_src2_reg[13]~128 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[13]~128 .shared_arith = "off";

dffeas \E_src2[13] (
	.clk(clk_clk),
	.d(\D_iw[19]~q ),
	.asdata(\D_src2_reg[13]~128_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[13]~q ),
	.prn(vcc));
defparam \E_src2[13] .is_wysiwyg = "true";
defparam \E_src2[13] .power_up = "low";

cyclonev_lcell_comb \Add17~9 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[7]~q ),
	.datae(gnd),
	.dataf(!\E_src1[7]~q ),
	.datag(gnd),
	.cin(\Add17~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~9_sumout ),
	.cout(\Add17~10 ),
	.shareout());
defparam \Add17~9 .extended_lut = "off";
defparam \Add17~9 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~9 .shared_arith = "off";

cyclonev_lcell_comb \Add17~1 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[8]~q ),
	.datae(gnd),
	.dataf(!\E_src1[8]~q ),
	.datag(gnd),
	.cin(\Add17~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~1_sumout ),
	.cout(\Add17~2 ),
	.shareout());
defparam \Add17~1 .extended_lut = "off";
defparam \Add17~1 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~1 .shared_arith = "off";

cyclonev_lcell_comb \Add17~5 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[9]~q ),
	.datae(gnd),
	.dataf(!\E_src1[9]~q ),
	.datag(gnd),
	.cin(\Add17~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~5_sumout ),
	.cout(\Add17~6 ),
	.shareout());
defparam \Add17~5 .extended_lut = "off";
defparam \Add17~5 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~5 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[9]~4 (
	.dataa(!\E_src2[9]~q ),
	.datab(!\E_src1[9]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[9]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[9]~4 .extended_lut = "off";
defparam \E_logic_result[9]~4 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[9]~4 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[9]~6 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[9]~4_combout ),
	.datad(!\E_extra_pc[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[9]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[9]~6 .extended_lut = "off";
defparam \E_alu_result[9]~6 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[9]~6 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[9] (
	.dataa(!\Add17~5_sumout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_alu_result[9]~6_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[9]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[9] .extended_lut = "off";
defparam \E_alu_result[9] .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \E_alu_result[9] .shared_arith = "off";

dffeas \M_alu_result[9] (
	.clk(clk_clk),
	.d(\E_alu_result[9]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[9]~q ),
	.prn(vcc));
defparam \M_alu_result[9] .is_wysiwyg = "true";
defparam \M_alu_result[9] .power_up = "low";

dffeas \A_inst_result[9] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[9] ),
	.asdata(\M_alu_result[9]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[9]~q ),
	.prn(vcc));
defparam \A_inst_result[9] .is_wysiwyg = "true";
defparam \A_inst_result[9] .power_up = "low";

dffeas A_ld_align_byte1_fill(
	.clk(clk_clk),
	.d(\M_ctrl_ld8~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ld_align_byte1_fill~q ),
	.prn(vcc));
defparam A_ld_align_byte1_fill.is_wysiwyg = "true";
defparam A_ld_align_byte1_fill.power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte1_data_aligned_nxt[1]~4 (
	.dataa(!\A_ld_align_sh16~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!\d_readdata_d1[25]~q ),
	.datae(!\d_readdata_d1[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte1_data_aligned_nxt[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte1_data_aligned_nxt[1]~4 .extended_lut = "off";
defparam \A_slow_ld_byte1_data_aligned_nxt[1]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_slow_ld_byte1_data_aligned_nxt[1]~4 .shared_arith = "off";

dffeas \A_slow_inst_result[9] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte1_data_aligned_nxt[1]~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[9]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[9] .is_wysiwyg = "true";
defparam \A_slow_inst_result[9] .power_up = "low";

cyclonev_lcell_comb A_data_ram_ld_align_fill_bit(
	.dataa(!\A_data_ram_ld_align_sign_bit~q ),
	.datab(!\A_ctrl_ld_signed~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_data_ram_ld_align_fill_bit~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_data_ram_ld_align_fill_bit.extended_lut = "off";
defparam A_data_ram_ld_align_fill_bit.lut_mask = 64'h7777777777777777;
defparam A_data_ram_ld_align_fill_bit.shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[11]~4 (
	.dataa(!\A_slow_inst_sel~q ),
	.datab(!\A_ld_align_sh16~q ),
	.datac(!\A_ld_align_byte1_fill~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[11]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[11]~4 .extended_lut = "off";
defparam \A_wr_data_unfiltered[11]~4 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \A_wr_data_unfiltered[11]~4 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[11]~5 (
	.dataa(!\A_slow_inst_sel~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[11]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[11]~5 .extended_lut = "off";
defparam \A_wr_data_unfiltered[11]~5 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_wr_data_unfiltered[11]~5 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[9]~14 (
	.dataa(!\A_inst_result[9]~q ),
	.datab(!\A_inst_result[25]~q ),
	.datac(!\A_slow_inst_result[9]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[11]~4_combout ),
	.dataf(!\A_wr_data_unfiltered[11]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[9]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[9]~14 .extended_lut = "off";
defparam \A_wr_data_unfiltered[9]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[9]~14 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[9]~12 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\A_mul_result[9]~q ),
	.datae(!\A_shift_rot_result[9]~q ),
	.dataf(!\A_wr_data_unfiltered[9]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[9]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[9]~12 .extended_lut = "off";
defparam \D_src2_reg[9]~12 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[9]~12 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[9]~96 (
	.dataa(!\M_alu_result[9]~q ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[5]~3_combout ),
	.datad(!\D_src2_reg[13]~8_combout ),
	.datae(!\W_wr_data[9]~q ),
	.dataf(!\D_src2_reg[9]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[9]~96_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[9]~96 .extended_lut = "off";
defparam \D_src2_reg[9]~96 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[9]~96 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[9]~112 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[9] ),
	.datad(!\D_src2_reg[9]~96_combout ),
	.datae(!\D_src2_reg[5]~2_combout ),
	.dataf(!\E_alu_result[9]~6_combout ),
	.datag(!\Add17~5_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[9]~112_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[9]~112 .extended_lut = "on";
defparam \D_src2_reg[9]~112 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[9]~112 .shared_arith = "off";

dffeas \E_src2[9] (
	.clk(clk_clk),
	.d(\D_iw[15]~q ),
	.asdata(\D_src2_reg[9]~112_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[9]~q ),
	.prn(vcc));
defparam \E_src2[9] .is_wysiwyg = "true";
defparam \E_src2[9] .power_up = "low";

cyclonev_lcell_comb \Add17~13 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[10]~q ),
	.datae(gnd),
	.dataf(!\E_src1[10]~q ),
	.datag(gnd),
	.cin(\Add17~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~13_sumout ),
	.cout(\Add17~14 ),
	.shareout());
defparam \Add17~13 .extended_lut = "off";
defparam \Add17~13 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~13 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[10]~3 (
	.dataa(!\E_src2[10]~q ),
	.datab(!\E_src1[10]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[10]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[10]~3 .extended_lut = "off";
defparam \E_logic_result[10]~3 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[10]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[10]~5 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[10]~3_combout ),
	.datad(!\E_extra_pc[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[10]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[10]~5 .extended_lut = "off";
defparam \E_alu_result[10]~5 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[10]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[10] (
	.dataa(!\Add17~13_sumout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_alu_result[10]~5_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[10]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[10] .extended_lut = "off";
defparam \E_alu_result[10] .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \E_alu_result[10] .shared_arith = "off";

dffeas \M_alu_result[10] (
	.clk(clk_clk),
	.d(\E_alu_result[10]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[10]~q ),
	.prn(vcc));
defparam \M_alu_result[10] .is_wysiwyg = "true";
defparam \M_alu_result[10] .power_up = "low";

dffeas \A_inst_result[10] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[10] ),
	.asdata(\M_alu_result[10]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[10]~q ),
	.prn(vcc));
defparam \A_inst_result[10] .is_wysiwyg = "true";
defparam \A_inst_result[10] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte1_data_aligned_nxt[2]~3 (
	.dataa(!\A_ld_align_sh16~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!\d_readdata_d1[26]~q ),
	.datae(!\d_readdata_d1[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte1_data_aligned_nxt[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte1_data_aligned_nxt[2]~3 .extended_lut = "off";
defparam \A_slow_ld_byte1_data_aligned_nxt[2]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_slow_ld_byte1_data_aligned_nxt[2]~3 .shared_arith = "off";

dffeas \A_slow_inst_result[10] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte1_data_aligned_nxt[2]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[10]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[10] .is_wysiwyg = "true";
defparam \A_slow_inst_result[10] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[10]~12 (
	.dataa(!\A_inst_result[10]~q ),
	.datab(!\A_inst_result[26]~q ),
	.datac(!\A_slow_inst_result[10]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[11]~4_combout ),
	.dataf(!\A_wr_data_unfiltered[11]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[10]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[10]~12 .extended_lut = "off";
defparam \A_wr_data_unfiltered[10]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[10]~12 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[10]~11 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\A_mul_result[10]~q ),
	.datae(!\A_shift_rot_result[10]~q ),
	.dataf(!\A_wr_data_unfiltered[10]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[10]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[10]~11 .extended_lut = "off";
defparam \D_src2_reg[10]~11 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[10]~11 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[10]~95 (
	.dataa(!\M_alu_result[10]~q ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[5]~3_combout ),
	.datad(!\D_src2_reg[13]~8_combout ),
	.datae(!\W_wr_data[10]~q ),
	.dataf(!\D_src2_reg[10]~11_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[10]~95_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[10]~95 .extended_lut = "off";
defparam \D_src2_reg[10]~95 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[10]~95 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[10]~116 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[10] ),
	.datad(!\D_src2_reg[10]~95_combout ),
	.datae(!\D_src2_reg[5]~2_combout ),
	.dataf(!\E_alu_result[10]~5_combout ),
	.datag(!\Add17~13_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[10]~116_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[10]~116 .extended_lut = "on";
defparam \D_src2_reg[10]~116 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[10]~116 .shared_arith = "off";

dffeas \E_src2[10] (
	.clk(clk_clk),
	.d(\D_iw[16]~q ),
	.asdata(\D_src2_reg[10]~116_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[10]~q ),
	.prn(vcc));
defparam \E_src2[10] .is_wysiwyg = "true";
defparam \E_src2[10] .power_up = "low";

cyclonev_lcell_comb \Add17~49 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[11]~q ),
	.datae(gnd),
	.dataf(!\E_src1[11]~q ),
	.datag(gnd),
	.cin(\Add17~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~49_sumout ),
	.cout(\Add17~50 ),
	.shareout());
defparam \Add17~49 .extended_lut = "off";
defparam \Add17~49 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~49 .shared_arith = "off";

cyclonev_lcell_comb \Add17~45 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[12]~q ),
	.datae(gnd),
	.dataf(!\E_src1[12]~q ),
	.datag(gnd),
	.cin(\Add17~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~45_sumout ),
	.cout(\Add17~46 ),
	.shareout());
defparam \Add17~45 .extended_lut = "off";
defparam \Add17~45 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~45 .shared_arith = "off";

cyclonev_lcell_comb \Add17~41 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[13]~q ),
	.datae(gnd),
	.dataf(!\E_src1[13]~q ),
	.datag(gnd),
	.cin(\Add17~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~41_sumout ),
	.cout(\Add17~42 ),
	.shareout());
defparam \Add17~41 .extended_lut = "off";
defparam \Add17~41 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~41 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[13] (
	.dataa(!\Add17~41_sumout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_alu_result[13]~2_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[13]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[13] .extended_lut = "off";
defparam \E_alu_result[13] .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \E_alu_result[13] .shared_arith = "off";

dffeas \M_alu_result[13] (
	.clk(clk_clk),
	.d(\E_alu_result[13]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[13]~q ),
	.prn(vcc));
defparam \M_alu_result[13] .is_wysiwyg = "true";
defparam \M_alu_result[13] .power_up = "low";

dffeas \A_inst_result[13] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[13] ),
	.asdata(\M_alu_result[13]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[13]~q ),
	.prn(vcc));
defparam \A_inst_result[13] .is_wysiwyg = "true";
defparam \A_inst_result[13] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte1_data_aligned_nxt[5]~0 (
	.dataa(!\A_ld_align_sh16~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!\d_readdata_d1[29]~q ),
	.datae(!\d_readdata_d1[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte1_data_aligned_nxt[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte1_data_aligned_nxt[5]~0 .extended_lut = "off";
defparam \A_slow_ld_byte1_data_aligned_nxt[5]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_slow_ld_byte1_data_aligned_nxt[5]~0 .shared_arith = "off";

dffeas \A_slow_inst_result[13] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte1_data_aligned_nxt[5]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[13]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[13] .is_wysiwyg = "true";
defparam \A_slow_inst_result[13] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[13]~6 (
	.dataa(!\A_inst_result[13]~q ),
	.datab(!\A_inst_result[29]~q ),
	.datac(!\A_slow_inst_result[13]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[11]~4_combout ),
	.dataf(!\A_wr_data_unfiltered[11]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[13]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[13]~6 .extended_lut = "off";
defparam \A_wr_data_unfiltered[13]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[13]~6 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[13]~7 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_mul_result[13]~q ),
	.datac(!\A_shift_rot_result[13]~q ),
	.datad(!\A_ctrl_shift_rot~q ),
	.datae(!\A_wr_data_unfiltered[13]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[13]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[13]~7 .extended_lut = "off";
defparam \A_wr_data_unfiltered[13]~7 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \A_wr_data_unfiltered[13]~7 .shared_arith = "off";

dffeas \W_wr_data[13] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[13]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[13]~q ),
	.prn(vcc));
defparam \W_wr_data[13] .is_wysiwyg = "true";
defparam \W_wr_data[13] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[13]~1 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[13] ),
	.datab(!\W_wr_data[13]~q ),
	.datac(!\M_alu_result[13]~q ),
	.datad(!\A_wr_data_unfiltered[13]~7_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[13]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[13]~1 .extended_lut = "off";
defparam \D_src1_reg[13]~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[13]~1 .shared_arith = "off";

dffeas \E_src1[13] (
	.clk(clk_clk),
	.d(\D_src1_reg[13]~1_combout ),
	.asdata(\E_alu_result[13]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[13]~q ),
	.prn(vcc));
defparam \E_src1[13] .is_wysiwyg = "true";
defparam \E_src1[13] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[13]~9 (
	.dataa(!\E_src1[13]~q ),
	.datab(!\E_src1[12]~q ),
	.datac(!\E_src1[11]~q ),
	.datad(!\E_src1[10]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[13]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[13]~9 .extended_lut = "off";
defparam \E_rot_step1[13]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[13]~9 .shared_arith = "off";

dffeas \M_rot_prestep2[13] (
	.clk(clk_clk),
	.d(\E_rot_step1[9]~8_combout ),
	.asdata(\E_rot_step1[13]~9_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[13]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[13] .is_wysiwyg = "true";
defparam \M_rot_prestep2[13] .power_up = "low";

cyclonev_lcell_comb \M_rot[5]~28 (
	.dataa(!\M_rot_prestep2[29]~q ),
	.datab(!\M_rot_prestep2[21]~q ),
	.datac(!\M_rot_prestep2[13]~q ),
	.datad(!\M_rot_prestep2[5]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~28 .extended_lut = "off";
defparam \M_rot[5]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~28 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~28 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[5]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[5]~28_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~28 .extended_lut = "off";
defparam \A_shift_rot_result~28 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~28 .shared_arith = "off";

dffeas \A_shift_rot_result[29] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~28_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[29]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[29] .is_wysiwyg = "true";
defparam \A_shift_rot_result[29] .power_up = "low";

dffeas \A_slow_inst_result[29] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[29]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[29]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[29] .is_wysiwyg = "true";
defparam \A_slow_inst_result[29] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[29]~59 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[29]~q ),
	.dataf(!\A_slow_inst_result[29]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[29]~59_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[29]~59 .extended_lut = "off";
defparam \A_wr_data_unfiltered[29]~59 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[29]~59 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[29]~60 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[29]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[29]~q ),
	.datae(!\A_wr_data_unfiltered[29]~59_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[29]~60_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[29]~60 .extended_lut = "off";
defparam \A_wr_data_unfiltered[29]~60 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[29]~60 .shared_arith = "off";

dffeas \W_wr_data[29] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[29]~60_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[29]~q ),
	.prn(vcc));
defparam \W_wr_data[29] .is_wysiwyg = "true";
defparam \W_wr_data[29] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[29]~13 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[29] ),
	.datab(!\W_wr_data[29]~q ),
	.datac(!\M_alu_result[29]~q ),
	.datad(!\A_wr_data_unfiltered[29]~60_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[29]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[29]~13 .extended_lut = "off";
defparam \D_src1_reg[29]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[29]~13 .shared_arith = "off";

dffeas \E_src1[29] (
	.clk(clk_clk),
	.d(\D_src1_reg[29]~13_combout ),
	.asdata(\E_alu_result[29]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[29]~q ),
	.prn(vcc));
defparam \E_src1[29] .is_wysiwyg = "true";
defparam \E_src1[29] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[29]~13 (
	.dataa(!\E_src1[29]~q ),
	.datab(!\E_src1[28]~q ),
	.datac(!\E_src1[27]~q ),
	.datad(!\E_src1[26]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[29]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[29]~13 .extended_lut = "off";
defparam \E_rot_step1[29]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[29]~13 .shared_arith = "off";

dffeas \M_rot_prestep2[1] (
	.clk(clk_clk),
	.d(\E_rot_step1[29]~13_combout ),
	.asdata(\E_rot_step1[1]~10_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[1]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[1] .is_wysiwyg = "true";
defparam \M_rot_prestep2[1] .power_up = "low";

dffeas \M_rot_prestep2[25] (
	.clk(clk_clk),
	.d(\E_rot_step1[21]~15_combout ),
	.asdata(\E_rot_step1[25]~12_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[25]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[25] .is_wysiwyg = "true";
defparam \M_rot_prestep2[25] .power_up = "low";

dffeas \M_rot_prestep2[17] (
	.clk(clk_clk),
	.d(\E_rot_step1[13]~9_combout ),
	.asdata(\E_rot_step1[17]~14_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[17]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[17] .is_wysiwyg = "true";
defparam \M_rot_prestep2[17] .power_up = "low";

cyclonev_lcell_comb \M_rot[1]~5 (
	.dataa(!\M_rot_prestep2[9]~q ),
	.datab(!\M_rot_prestep2[1]~q ),
	.datac(!\M_rot_prestep2[25]~q ),
	.datad(!\M_rot_prestep2[17]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~5 .extended_lut = "off";
defparam \M_rot[1]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~5 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~5 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_sel_fill1~q ),
	.datad(!\M_rot_mask[1]~q ),
	.datae(!\M_rot[1]~5_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~5 .extended_lut = "off";
defparam \A_shift_rot_result~5 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~5 .shared_arith = "off";

dffeas \A_shift_rot_result[9] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[9]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[9] .is_wysiwyg = "true";
defparam \A_shift_rot_result[9] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[9]~15 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[9]~q ),
	.datad(!\A_shift_rot_result[9]~q ),
	.datae(!\A_wr_data_unfiltered[9]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[9]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[9]~15 .extended_lut = "off";
defparam \A_wr_data_unfiltered[9]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[9]~15 .shared_arith = "off";

dffeas \W_wr_data[9] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[9]~15_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[9]~q ),
	.prn(vcc));
defparam \W_wr_data[9] .is_wysiwyg = "true";
defparam \W_wr_data[9] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[9]~5 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[9] ),
	.datab(!\W_wr_data[9]~q ),
	.datac(!\M_alu_result[9]~q ),
	.datad(!\A_wr_data_unfiltered[9]~15_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[9]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[9]~5 .extended_lut = "off";
defparam \D_src1_reg[9]~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[9]~5 .shared_arith = "off";

dffeas \E_src1[9] (
	.clk(clk_clk),
	.d(\D_src1_reg[9]~5_combout ),
	.asdata(\E_alu_result[9]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[9]~q ),
	.prn(vcc));
defparam \E_src1[9] .is_wysiwyg = "true";
defparam \E_src1[9] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[11]~25 (
	.dataa(!\E_src1[11]~q ),
	.datab(!\E_src1[10]~q ),
	.datac(!\E_src1[9]~q ),
	.datad(!\E_src1[8]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[11]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[11]~25 .extended_lut = "off";
defparam \E_rot_step1[11]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[11]~25 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[15]~30 (
	.dataa(!\E_src1[15]~q ),
	.datab(!\E_src1[14]~q ),
	.datac(!\E_src1[13]~q ),
	.datad(!\E_src1[12]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[15]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[15]~30 .extended_lut = "off";
defparam \E_rot_step1[15]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[15]~30 .shared_arith = "off";

dffeas \M_rot_prestep2[15] (
	.clk(clk_clk),
	.d(\E_rot_step1[11]~25_combout ),
	.asdata(\E_rot_step1[15]~30_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[15]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[15] .is_wysiwyg = "true";
defparam \M_rot_prestep2[15] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[3]~27 (
	.dataa(!\E_src1[3]~q ),
	.datab(!\E_src1[2]~q ),
	.datac(!\E_src1[1]~q ),
	.datad(!\E_src1[0]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[3]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[3]~27 .extended_lut = "off";
defparam \E_rot_step1[3]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[3]~27 .shared_arith = "off";

dffeas \M_rot_prestep2[7] (
	.clk(clk_clk),
	.d(\E_rot_step1[3]~27_combout ),
	.asdata(\E_rot_step1[7]~24_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[7]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[7] .is_wysiwyg = "true";
defparam \M_rot_prestep2[7] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[27]~29 (
	.dataa(!\E_src1[27]~q ),
	.datab(!\E_src1[26]~q ),
	.datac(!\E_src1[25]~q ),
	.datad(!\E_src1[24]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[27]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[27]~29 .extended_lut = "off";
defparam \E_rot_step1[27]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[27]~29 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[31]~26 (
	.dataa(!\E_src1[31]~q ),
	.datab(!\E_src1[30]~q ),
	.datac(!\E_src1[29]~q ),
	.datad(!\E_src1[28]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[31]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[31]~26 .extended_lut = "off";
defparam \E_rot_step1[31]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[31]~26 .shared_arith = "off";

dffeas \M_rot_prestep2[31] (
	.clk(clk_clk),
	.d(\E_rot_step1[27]~29_combout ),
	.asdata(\E_rot_step1[31]~26_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[31]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[31] .is_wysiwyg = "true";
defparam \M_rot_prestep2[31] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[19]~31 (
	.dataa(!\E_src1[19]~q ),
	.datab(!\E_src1[18]~q ),
	.datac(!\E_src1[17]~q ),
	.datad(!\E_src1[16]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[19]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[19]~31 .extended_lut = "off";
defparam \E_rot_step1[19]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[19]~31 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[23]~28 (
	.dataa(!\E_src1[23]~q ),
	.datab(!\E_src1[22]~q ),
	.datac(!\E_src1[21]~q ),
	.datad(!\E_src1[20]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[23]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[23]~28 .extended_lut = "off";
defparam \E_rot_step1[23]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[23]~28 .shared_arith = "off";

dffeas \M_rot_prestep2[23] (
	.clk(clk_clk),
	.d(\E_rot_step1[19]~31_combout ),
	.asdata(\E_rot_step1[23]~28_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[23]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[23] .is_wysiwyg = "true";
defparam \M_rot_prestep2[23] .power_up = "low";

cyclonev_lcell_comb \M_rot[7]~25 (
	.dataa(!\M_rot_prestep2[15]~q ),
	.datab(!\M_rot_prestep2[7]~q ),
	.datac(!\M_rot_prestep2[31]~q ),
	.datad(!\M_rot_prestep2[23]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~25 .extended_lut = "off";
defparam \M_rot[7]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~25 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~25 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_sel_fill1~q ),
	.datad(!\M_rot_mask[7]~q ),
	.datae(!\M_rot[7]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~25 .extended_lut = "off";
defparam \A_shift_rot_result~25 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~25 .shared_arith = "off";

dffeas \A_shift_rot_result[15] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~25_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[15]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[15] .is_wysiwyg = "true";
defparam \A_shift_rot_result[15] .power_up = "low";

dffeas \A_inst_result[15] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.asdata(\M_alu_result[15]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[15]~q ),
	.prn(vcc));
defparam \A_inst_result[15] .is_wysiwyg = "true";
defparam \A_inst_result[15] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte1_data_aligned_nxt[7]~6 (
	.dataa(!\A_ld_align_sh16~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(!\d_readdata_d1[15]~q ),
	.datad(!\d_readdata_d1[31]~q ),
	.datae(!\A_slow_ld_data_fill_bit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte1_data_aligned_nxt[7]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte1_data_aligned_nxt[7]~6 .extended_lut = "off";
defparam \A_slow_ld_byte1_data_aligned_nxt[7]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_slow_ld_byte1_data_aligned_nxt[7]~6 .shared_arith = "off";

dffeas \A_slow_inst_result[15] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte1_data_aligned_nxt[7]~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[15]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[15] .is_wysiwyg = "true";
defparam \A_slow_inst_result[15] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[15]~55 (
	.dataa(!\A_inst_result[15]~q ),
	.datab(!\A_inst_result[31]~q ),
	.datac(!\A_slow_inst_result[15]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[11]~4_combout ),
	.dataf(!\A_wr_data_unfiltered[11]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[15]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[15]~55 .extended_lut = "off";
defparam \A_wr_data_unfiltered[15]~55 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[15]~55 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[15]~67 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[15]~q ),
	.datad(!\A_shift_rot_result[15]~q ),
	.datae(!\A_wr_data_unfiltered[15]~55_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[15]~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[15]~67 .extended_lut = "off";
defparam \A_wr_data_unfiltered[15]~67 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[15]~67 .shared_arith = "off";

dffeas \W_wr_data[15] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[15]~67_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[15]~q ),
	.prn(vcc));
defparam \W_wr_data[15] .is_wysiwyg = "true";
defparam \W_wr_data[15] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[15]~23 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[15] ),
	.datab(!\W_wr_data[15]~q ),
	.datac(!\M_alu_result[15]~q ),
	.datad(!\A_wr_data_unfiltered[15]~67_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[15]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[15]~23 .extended_lut = "off";
defparam \D_src1_reg[15]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[15]~23 .shared_arith = "off";

dffeas \E_src1[15] (
	.clk(clk_clk),
	.d(\D_src1_reg[15]~23_combout ),
	.asdata(\E_alu_result[15]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[15]~q ),
	.prn(vcc));
defparam \E_src1[15] .is_wysiwyg = "true";
defparam \E_src1[15] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[15]~11 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[15]~q ),
	.datad(!\E_src1[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[15]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[15]~11 .extended_lut = "off";
defparam \E_logic_result[15]~11 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[15]~11 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~25 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[15]~11_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~25 .extended_lut = "off";
defparam \E_alu_result~25 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~25 .shared_arith = "off";

cyclonev_lcell_comb \Add17~125 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[14]~q ),
	.datae(gnd),
	.dataf(!\E_src1[14]~q ),
	.datag(gnd),
	.cin(\Add17~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~125_sumout ),
	.cout(\Add17~126 ),
	.shareout());
defparam \Add17~125 .extended_lut = "off";
defparam \Add17~125 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~125 .shared_arith = "off";

cyclonev_lcell_comb \Add17~117 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[15]~q ),
	.datae(gnd),
	.dataf(!\E_src1[15]~q ),
	.datag(gnd),
	.cin(\Add17~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~117_sumout ),
	.cout(\Add17~118 ),
	.shareout());
defparam \Add17~117 .extended_lut = "off";
defparam \Add17~117 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~117 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[15] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~25_combout ),
	.datac(!\Add17~117_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[15]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[15] .extended_lut = "off";
defparam \E_alu_result[15] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[15] .shared_arith = "off";

dffeas \M_alu_result[15] (
	.clk(clk_clk),
	.d(\E_alu_result[15]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[15]~q ),
	.prn(vcc));
defparam \M_alu_result[15] .is_wysiwyg = "true";
defparam \M_alu_result[15] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[15]~51 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\A_mul_result[15]~q ),
	.datae(!\A_shift_rot_result[15]~q ),
	.dataf(!\A_wr_data_unfiltered[15]~55_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[15]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[15]~51 .extended_lut = "off";
defparam \D_src2_reg[15]~51 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[15]~51 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[15]~98 (
	.dataa(!\D_src2_reg[5]~4_combout ),
	.datab(!\M_alu_result[15]~q ),
	.datac(!\D_src2_reg[5]~3_combout ),
	.datad(!\D_src2_reg[13]~8_combout ),
	.datae(!\W_wr_data[15]~q ),
	.dataf(!\D_src2_reg[15]~51_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[15]~98_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[15]~98 .extended_lut = "off";
defparam \D_src2_reg[15]~98 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \D_src2_reg[15]~98 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[15]~104 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[15] ),
	.datad(!\D_src2_reg[15]~98_combout ),
	.datae(!\D_src2_reg[5]~2_combout ),
	.dataf(!\Add17~117_sumout ),
	.datag(!\E_alu_result~25_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[15]~104_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[15]~104 .extended_lut = "on";
defparam \D_src2_reg[15]~104 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[15]~104 .shared_arith = "off";

dffeas \E_src2[15] (
	.clk(clk_clk),
	.d(\D_iw[21]~q ),
	.asdata(\D_src2_reg[15]~104_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[15]~q ),
	.prn(vcc));
defparam \E_src2[15] .is_wysiwyg = "true";
defparam \E_src2[15] .power_up = "low";

cyclonev_lcell_comb \Add17~93 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[16]~q ),
	.datae(gnd),
	.dataf(!\E_src1[16]~q ),
	.datag(gnd),
	.cin(\Add17~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~93_sumout ),
	.cout(\Add17~94 ),
	.shareout());
defparam \Add17~93 .extended_lut = "off";
defparam \Add17~93 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~93 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[16] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~19_combout ),
	.datac(!\Add17~93_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[16]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[16] .extended_lut = "off";
defparam \E_alu_result[16] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[16] .shared_arith = "off";

dffeas \M_alu_result[16] (
	.clk(clk_clk),
	.d(\E_alu_result[16]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[16]~q ),
	.prn(vcc));
defparam \M_alu_result[16] .is_wysiwyg = "true";
defparam \M_alu_result[16] .power_up = "low";

dffeas \A_inst_result[16] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[16] ),
	.asdata(\M_alu_result[16]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[16]~q ),
	.prn(vcc));
defparam \A_inst_result[16] .is_wysiwyg = "true";
defparam \A_inst_result[16] .power_up = "low";

cyclonev_lcell_comb \E_rot_pass2~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(!\E_ctrl_shift_rot_left~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass2~0 .extended_lut = "off";
defparam \E_rot_pass2~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \E_rot_pass2~0 .shared_arith = "off";

dffeas M_rot_pass2(
	.clk(clk_clk),
	.d(\E_rot_pass2~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_pass2~q ),
	.prn(vcc));
defparam M_rot_pass2.is_wysiwyg = "true";
defparam M_rot_pass2.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill2~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_right~q ),
	.datad(!\E_ctrl_shift_rot_left~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill2~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill2~0 .extended_lut = "off";
defparam \E_rot_sel_fill2~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_sel_fill2~0 .shared_arith = "off";

dffeas M_rot_sel_fill2(
	.clk(clk_clk),
	.d(\E_rot_sel_fill2~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_sel_fill2~q ),
	.prn(vcc));
defparam M_rot_sel_fill2.is_wysiwyg = "true";
defparam M_rot_sel_fill2.power_up = "low";

cyclonev_lcell_comb \E_rot_step1[12]~17 (
	.dataa(!\E_src1[12]~q ),
	.datab(!\E_src1[11]~q ),
	.datac(!\E_src1[10]~q ),
	.datad(!\E_src1[9]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[12]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[12]~17 .extended_lut = "off";
defparam \E_rot_step1[12]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[12]~17 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[16]~22 (
	.dataa(!\E_src1[16]~q ),
	.datab(!\E_src1[15]~q ),
	.datac(!\E_src1[14]~q ),
	.datad(!\E_src1[13]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[16]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[16]~22 .extended_lut = "off";
defparam \E_rot_step1[16]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[16]~22 .shared_arith = "off";

dffeas \M_rot_prestep2[16] (
	.clk(clk_clk),
	.d(\E_rot_step1[12]~17_combout ),
	.asdata(\E_rot_step1[16]~22_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[16]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[16] .is_wysiwyg = "true";
defparam \M_rot_prestep2[16] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[20]~23 (
	.dataa(!\E_src1[20]~q ),
	.datab(!\E_src1[19]~q ),
	.datac(!\E_src1[18]~q ),
	.datad(!\E_src1[17]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[20]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[20]~23 .extended_lut = "off";
defparam \E_rot_step1[20]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[20]~23 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_step1[24]~20 (
	.dataa(!\E_src1[24]~q ),
	.datab(!\E_src1[23]~q ),
	.datac(!\E_src1[22]~q ),
	.datad(!\E_src1[21]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[24]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[24]~20 .extended_lut = "off";
defparam \E_rot_step1[24]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[24]~20 .shared_arith = "off";

dffeas \M_rot_prestep2[24] (
	.clk(clk_clk),
	.d(\E_rot_step1[20]~23_combout ),
	.asdata(\E_rot_step1[24]~20_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[24]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[24] .is_wysiwyg = "true";
defparam \M_rot_prestep2[24] .power_up = "low";

cyclonev_lcell_comb \M_rot[0]~19 (
	.dataa(!\M_rot_prestep2[16]~q ),
	.datab(!\M_rot_prestep2[8]~q ),
	.datac(!\M_rot_prestep2[0]~q ),
	.datad(!\M_rot_prestep2[24]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~19 .extended_lut = "off";
defparam \M_rot[0]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~19 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~19 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[0]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[0]~19_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~19 .extended_lut = "off";
defparam \A_shift_rot_result~19 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~19 .shared_arith = "off";

dffeas \A_shift_rot_result[16] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~19_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[16]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[16] .is_wysiwyg = "true";
defparam \A_shift_rot_result[16] .power_up = "low";

dffeas \A_slow_inst_result[16] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[16]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[16]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[16] .is_wysiwyg = "true";
defparam \A_slow_inst_result[16] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[16]~43 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[16]~q ),
	.dataf(!\A_slow_inst_result[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[16]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[16]~43 .extended_lut = "off";
defparam \A_wr_data_unfiltered[16]~43 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[16]~43 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[16]~44 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[16]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[16]~q ),
	.datae(!\A_wr_data_unfiltered[16]~43_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[16]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[16]~44 .extended_lut = "off";
defparam \A_wr_data_unfiltered[16]~44 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[16]~44 .shared_arith = "off";

dffeas \W_wr_data[16] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[16]~44_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[16]~q ),
	.prn(vcc));
defparam \W_wr_data[16] .is_wysiwyg = "true";
defparam \W_wr_data[16] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[16]~39 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\W_wr_data[16]~q ),
	.datad(!\A_wr_data_unfiltered[16]~44_combout ),
	.datae(!\M_alu_result[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[16]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[16]~39 .extended_lut = "off";
defparam \D_src2_reg[16]~39 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[16]~39 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[16]~32 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\D_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\D_ctrl_unsigned_lo_imm16~q ),
	.dataf(!\D_iw[6]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[16]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[16]~32 .extended_lut = "off";
defparam \D_src2[16]~32 .lut_mask = 64'hEDFFDEFFFFFFFFFF;
defparam \D_src2[16]~32 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[16]~33 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_alu_result~19_combout ),
	.datac(!\Add17~93_sumout ),
	.datad(!\D_src2[16]~32_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[16]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[16]~33 .extended_lut = "off";
defparam \D_src2[16]~33 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \D_src2[16]~33 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[16]~9 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_ctrl_src2_choose_imm~q ),
	.datad(!\D_src2_reg[16]~39_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(!\D_src2[16]~33_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[16]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[16]~9 .extended_lut = "off";
defparam \D_src2[16]~9 .lut_mask = 64'hFFFFFFFF96FFFFFF;
defparam \D_src2[16]~9 .shared_arith = "off";

dffeas \E_src2[16] (
	.clk(clk_clk),
	.d(\D_src2[16]~9_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[16]~q ),
	.prn(vcc));
defparam \E_src2[16] .is_wysiwyg = "true";
defparam \E_src2[16] .power_up = "low";

cyclonev_lcell_comb \Add17~85 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[17]~q ),
	.datae(gnd),
	.dataf(!\E_src1[17]~q ),
	.datag(gnd),
	.cin(\Add17~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~85_sumout ),
	.cout(\Add17~86 ),
	.shareout());
defparam \Add17~85 .extended_lut = "off";
defparam \Add17~85 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~85 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[17] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~17_combout ),
	.datac(!\Add17~85_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[17]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[17] .extended_lut = "off";
defparam \E_alu_result[17] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[17] .shared_arith = "off";

dffeas \M_alu_result[17] (
	.clk(clk_clk),
	.d(\E_alu_result[17]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[17]~q ),
	.prn(vcc));
defparam \M_alu_result[17] .is_wysiwyg = "true";
defparam \M_alu_result[17] .power_up = "low";

dffeas \A_inst_result[17] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[17] ),
	.asdata(\M_alu_result[17]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[17]~q ),
	.prn(vcc));
defparam \A_inst_result[17] .is_wysiwyg = "true";
defparam \A_inst_result[17] .power_up = "low";

cyclonev_lcell_comb \M_rot[1]~17 (
	.dataa(!\M_rot_prestep2[17]~q ),
	.datab(!\M_rot_prestep2[9]~q ),
	.datac(!\M_rot_prestep2[1]~q ),
	.datad(!\M_rot_prestep2[25]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~17 .extended_lut = "off";
defparam \M_rot[1]~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~17 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~17 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[1]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[1]~17_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~17 .extended_lut = "off";
defparam \A_shift_rot_result~17 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~17 .shared_arith = "off";

dffeas \A_shift_rot_result[17] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~17_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[17]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[17] .is_wysiwyg = "true";
defparam \A_shift_rot_result[17] .power_up = "low";

dffeas \A_slow_inst_result[17] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[17]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[17]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[17] .is_wysiwyg = "true";
defparam \A_slow_inst_result[17] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[17]~39 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[17]~q ),
	.dataf(!\A_slow_inst_result[17]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[17]~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[17]~39 .extended_lut = "off";
defparam \A_wr_data_unfiltered[17]~39 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[17]~39 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[17]~40 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[17]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[17]~q ),
	.datae(!\A_wr_data_unfiltered[17]~39_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[17]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[17]~40 .extended_lut = "off";
defparam \A_wr_data_unfiltered[17]~40 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[17]~40 .shared_arith = "off";

dffeas \W_wr_data[17] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[17]~40_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[17]~q ),
	.prn(vcc));
defparam \W_wr_data[17] .is_wysiwyg = "true";
defparam \W_wr_data[17] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[17]~35 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\W_wr_data[17]~q ),
	.datad(!\A_wr_data_unfiltered[17]~40_combout ),
	.datae(!\M_alu_result[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[17]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[17]~35 .extended_lut = "off";
defparam \D_src2_reg[17]~35 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[17]~35 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[17]~30 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\D_ctrl_hi_imm16~q ),
	.datad(!\D_iw[21]~q ),
	.datae(!\D_ctrl_unsigned_lo_imm16~q ),
	.dataf(!\D_iw[7]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[17]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[17]~30 .extended_lut = "off";
defparam \D_src2[17]~30 .lut_mask = 64'hEDFFDEFFFFFFFFFF;
defparam \D_src2[17]~30 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[17]~31 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\E_alu_result~17_combout ),
	.datac(!\Add17~85_sumout ),
	.datad(!\D_src2[17]~30_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[17]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[17]~31 .extended_lut = "off";
defparam \D_src2[17]~31 .lut_mask = 64'hFFD8FFD8FFD8FFD8;
defparam \D_src2[17]~31 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[17]~8 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_ctrl_src2_choose_imm~q ),
	.datad(!\D_src2_reg[17]~35_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(!\D_src2[17]~31_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[17]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[17]~8 .extended_lut = "off";
defparam \D_src2[17]~8 .lut_mask = 64'hFFFFFFFF96FFFFFF;
defparam \D_src2[17]~8 .shared_arith = "off";

dffeas \E_src2[17] (
	.clk(clk_clk),
	.d(\D_src2[17]~8_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[17]~q ),
	.prn(vcc));
defparam \E_src2[17] .is_wysiwyg = "true";
defparam \E_src2[17] .power_up = "low";

cyclonev_lcell_comb \Add17~109 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[18]~q ),
	.datae(gnd),
	.dataf(!\E_src1[18]~q ),
	.datag(gnd),
	.cin(\Add17~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~109_sumout ),
	.cout(\Add17~110 ),
	.shareout());
defparam \Add17~109 .extended_lut = "off";
defparam \Add17~109 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~109 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[18] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~23_combout ),
	.datac(!\Add17~109_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[18]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[18] .extended_lut = "off";
defparam \E_alu_result[18] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[18] .shared_arith = "off";

dffeas \M_alu_result[18] (
	.clk(clk_clk),
	.d(\E_alu_result[18]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[18]~q ),
	.prn(vcc));
defparam \M_alu_result[18] .is_wysiwyg = "true";
defparam \M_alu_result[18] .power_up = "low";

dffeas \A_inst_result[18] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[18] ),
	.asdata(\M_alu_result[18]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[18]~q ),
	.prn(vcc));
defparam \A_inst_result[18] .is_wysiwyg = "true";
defparam \A_inst_result[18] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[14]~4 (
	.dataa(!\E_src1[14]~q ),
	.datab(!\E_src1[13]~q ),
	.datac(!\E_src1[12]~q ),
	.datad(!\E_src1[11]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[14]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[14]~4 .extended_lut = "off";
defparam \E_rot_step1[14]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[14]~4 .shared_arith = "off";

dffeas \M_rot_prestep2[18] (
	.clk(clk_clk),
	.d(\E_rot_step1[14]~4_combout ),
	.asdata(\E_rot_step1[18]~5_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[18]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[18] .is_wysiwyg = "true";
defparam \M_rot_prestep2[18] .power_up = "low";

dffeas \M_rot_prestep2[2] (
	.clk(clk_clk),
	.d(\E_rot_step1[30]~0_combout ),
	.asdata(\E_rot_step1[2]~1_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[2]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[2] .is_wysiwyg = "true";
defparam \M_rot_prestep2[2] .power_up = "low";

dffeas \M_rot_prestep2[26] (
	.clk(clk_clk),
	.d(\E_rot_step1[22]~2_combout ),
	.asdata(\E_rot_step1[26]~3_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[26]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[26] .is_wysiwyg = "true";
defparam \M_rot_prestep2[26] .power_up = "low";

cyclonev_lcell_comb \M_rot[2]~23 (
	.dataa(!\M_rot_prestep2[18]~q ),
	.datab(!\M_rot_prestep2[10]~q ),
	.datac(!\M_rot_prestep2[2]~q ),
	.datad(!\M_rot_prestep2[26]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~23 .extended_lut = "off";
defparam \M_rot[2]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~23 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~23 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[2]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[2]~23_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~23 .extended_lut = "off";
defparam \A_shift_rot_result~23 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~23 .shared_arith = "off";

dffeas \A_shift_rot_result[18] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~23_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[18]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[18] .is_wysiwyg = "true";
defparam \A_shift_rot_result[18] .power_up = "low";

dffeas \A_slow_inst_result[18] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[18]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[18]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[18] .is_wysiwyg = "true";
defparam \A_slow_inst_result[18] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[18]~51 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[18]~q ),
	.dataf(!\A_slow_inst_result[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[18]~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[18]~51 .extended_lut = "off";
defparam \A_wr_data_unfiltered[18]~51 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[18]~51 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[18]~52 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[18]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[18]~q ),
	.datae(!\A_wr_data_unfiltered[18]~51_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[18]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[18]~52 .extended_lut = "off";
defparam \A_wr_data_unfiltered[18]~52 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[18]~52 .shared_arith = "off";

dffeas \W_wr_data[18] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[18]~52_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[18]~q ),
	.prn(vcc));
defparam \W_wr_data[18] .is_wysiwyg = "true";
defparam \W_wr_data[18] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[18]~19 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[18] ),
	.datab(!\W_wr_data[18]~q ),
	.datac(!\M_alu_result[18]~q ),
	.datad(!\A_wr_data_unfiltered[18]~52_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[18]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[18]~19 .extended_lut = "off";
defparam \D_src1_reg[18]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[18]~19 .shared_arith = "off";

dffeas \E_src1[18] (
	.clk(clk_clk),
	.d(\D_src1_reg[18]~19_combout ),
	.asdata(\E_alu_result[18]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[18]~q ),
	.prn(vcc));
defparam \E_src1[18] .is_wysiwyg = "true";
defparam \E_src1[18] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~23 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[18]~q ),
	.datae(!\E_src1[18]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~23 .extended_lut = "off";
defparam \E_alu_result~23 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~23 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[18]~65 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~23_combout ),
	.datad(!\Add17~109_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[18]~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[18]~65 .extended_lut = "off";
defparam \D_src2_reg[18]~65 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[18]~65 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[18]~47 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[18]~q ),
	.datae(!\A_wr_data_unfiltered[18]~52_combout ),
	.dataf(!\M_alu_result[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[18]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[18]~47 .extended_lut = "off";
defparam \D_src2_reg[18]~47 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[18]~47 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[18]~12 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[8]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[18]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[18]~12 .extended_lut = "off";
defparam \D_src2[18]~12 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \D_src2[18]~12 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[18]~13 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[18]~65_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.datae(!\D_src2_reg[18]~47_combout ),
	.dataf(!\D_src2[18]~12_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[18]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[18]~13 .extended_lut = "off";
defparam \D_src2[18]~13 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[18]~13 .shared_arith = "off";

dffeas \E_src2[18] (
	.clk(clk_clk),
	.d(\D_src2[18]~13_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[18]~q ),
	.prn(vcc));
defparam \E_src2[18] .is_wysiwyg = "true";
defparam \E_src2[18] .power_up = "low";

cyclonev_lcell_comb \Add17~101 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[19]~q ),
	.datae(gnd),
	.dataf(!\E_src1[19]~q ),
	.datag(gnd),
	.cin(\Add17~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~101_sumout ),
	.cout(\Add17~102 ),
	.shareout());
defparam \Add17~101 .extended_lut = "off";
defparam \Add17~101 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~101 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[19] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~21_combout ),
	.datac(!\Add17~101_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[19]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[19] .extended_lut = "off";
defparam \E_alu_result[19] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[19] .shared_arith = "off";

dffeas \M_alu_result[19] (
	.clk(clk_clk),
	.d(\E_alu_result[19]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[19]~q ),
	.prn(vcc));
defparam \M_alu_result[19] .is_wysiwyg = "true";
defparam \M_alu_result[19] .power_up = "low";

dffeas \A_inst_result[19] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[19] ),
	.asdata(\M_alu_result[19]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[19]~q ),
	.prn(vcc));
defparam \A_inst_result[19] .is_wysiwyg = "true";
defparam \A_inst_result[19] .power_up = "low";

dffeas \M_rot_prestep2[19] (
	.clk(clk_clk),
	.d(\E_rot_step1[15]~30_combout ),
	.asdata(\E_rot_step1[19]~31_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[19]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[19] .is_wysiwyg = "true";
defparam \M_rot_prestep2[19] .power_up = "low";

dffeas \M_rot_prestep2[3] (
	.clk(clk_clk),
	.d(\E_rot_step1[31]~26_combout ),
	.asdata(\E_rot_step1[3]~27_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[3]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[3] .is_wysiwyg = "true";
defparam \M_rot_prestep2[3] .power_up = "low";

dffeas \M_rot_prestep2[27] (
	.clk(clk_clk),
	.d(\E_rot_step1[23]~28_combout ),
	.asdata(\E_rot_step1[27]~29_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[27]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[27] .is_wysiwyg = "true";
defparam \M_rot_prestep2[27] .power_up = "low";

cyclonev_lcell_comb \M_rot[3]~21 (
	.dataa(!\M_rot_prestep2[19]~q ),
	.datab(!\M_rot_prestep2[11]~q ),
	.datac(!\M_rot_prestep2[3]~q ),
	.datad(!\M_rot_prestep2[27]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~21 .extended_lut = "off";
defparam \M_rot[3]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~21 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~21 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[3]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[3]~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~21 .extended_lut = "off";
defparam \A_shift_rot_result~21 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~21 .shared_arith = "off";

dffeas \A_shift_rot_result[19] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~21_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[19]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[19] .is_wysiwyg = "true";
defparam \A_shift_rot_result[19] .power_up = "low";

dffeas \A_slow_inst_result[19] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[19]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[19]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[19] .is_wysiwyg = "true";
defparam \A_slow_inst_result[19] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[19]~47 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[19]~q ),
	.dataf(!\A_slow_inst_result[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[19]~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[19]~47 .extended_lut = "off";
defparam \A_wr_data_unfiltered[19]~47 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[19]~47 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[19]~48 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[19]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[19]~q ),
	.datae(!\A_wr_data_unfiltered[19]~47_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[19]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[19]~48 .extended_lut = "off";
defparam \A_wr_data_unfiltered[19]~48 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[19]~48 .shared_arith = "off";

dffeas \W_wr_data[19] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[19]~48_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[19]~q ),
	.prn(vcc));
defparam \W_wr_data[19] .is_wysiwyg = "true";
defparam \W_wr_data[19] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[19]~21 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[19] ),
	.datab(!\W_wr_data[19]~q ),
	.datac(!\M_alu_result[19]~q ),
	.datad(!\A_wr_data_unfiltered[19]~48_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[19]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[19]~21 .extended_lut = "off";
defparam \D_src1_reg[19]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[19]~21 .shared_arith = "off";

dffeas \E_src1[19] (
	.clk(clk_clk),
	.d(\D_src1_reg[19]~21_combout ),
	.asdata(\E_alu_result[19]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[19]~q ),
	.prn(vcc));
defparam \E_src1[19] .is_wysiwyg = "true";
defparam \E_src1[19] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~21 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[19]~q ),
	.datae(!\E_src1[19]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~21 .extended_lut = "off";
defparam \E_alu_result~21 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~21 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[19]~67 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~21_combout ),
	.datad(!\Add17~101_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[19]~67_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[19]~67 .extended_lut = "off";
defparam \D_src2_reg[19]~67 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[19]~67 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[19]~43 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[19]~q ),
	.datae(!\A_wr_data_unfiltered[19]~48_combout ),
	.dataf(!\M_alu_result[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[19]~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[19]~43 .extended_lut = "off";
defparam \D_src2_reg[19]~43 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[19]~43 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[19]~16 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[9]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[19]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[19]~16 .extended_lut = "off";
defparam \D_src2[19]~16 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \D_src2[19]~16 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[19]~17 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[19]~67_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.datae(!\D_src2_reg[19]~43_combout ),
	.dataf(!\D_src2[19]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[19]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[19]~17 .extended_lut = "off";
defparam \D_src2[19]~17 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[19]~17 .shared_arith = "off";

dffeas \E_src2[19] (
	.clk(clk_clk),
	.d(\D_src2[19]~17_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[19]~q ),
	.prn(vcc));
defparam \E_src2[19] .is_wysiwyg = "true";
defparam \E_src2[19] .power_up = "low";

cyclonev_lcell_comb \Add17~77 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[20]~q ),
	.datae(gnd),
	.dataf(!\E_src1[20]~q ),
	.datag(gnd),
	.cin(\Add17~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~77_sumout ),
	.cout(\Add17~78 ),
	.shareout());
defparam \Add17~77 .extended_lut = "off";
defparam \Add17~77 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~77 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[20] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~15_combout ),
	.datac(!\Add17~77_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[20]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[20] .extended_lut = "off";
defparam \E_alu_result[20] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[20] .shared_arith = "off";

dffeas \M_alu_result[20] (
	.clk(clk_clk),
	.d(\E_alu_result[20]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[20]~q ),
	.prn(vcc));
defparam \M_alu_result[20] .is_wysiwyg = "true";
defparam \M_alu_result[20] .power_up = "low";

dffeas \A_inst_result[20] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[20] ),
	.asdata(\M_alu_result[20]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[20]~q ),
	.prn(vcc));
defparam \A_inst_result[20] .is_wysiwyg = "true";
defparam \A_inst_result[20] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[4]~2 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[4]~2 .extended_lut = "off";
defparam \E_rot_mask[4]~2 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_rot_mask[4]~2 .shared_arith = "off";

dffeas \M_rot_mask[4] (
	.clk(clk_clk),
	.d(\E_rot_mask[4]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[4]~q ),
	.prn(vcc));
defparam \M_rot_mask[4] .is_wysiwyg = "true";
defparam \M_rot_mask[4] .power_up = "low";

dffeas \M_rot_prestep2[20] (
	.clk(clk_clk),
	.d(\E_rot_step1[16]~22_combout ),
	.asdata(\E_rot_step1[20]~23_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[20]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[20] .is_wysiwyg = "true";
defparam \M_rot_prestep2[20] .power_up = "low";

dffeas \M_rot_prestep2[12] (
	.clk(clk_clk),
	.d(\E_rot_step1[8]~16_combout ),
	.asdata(\E_rot_step1[12]~17_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[12]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[12] .is_wysiwyg = "true";
defparam \M_rot_prestep2[12] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[0]~18 (
	.dataa(!\E_src1[0]~q ),
	.datab(!\E_src1[31]~q ),
	.datac(!\E_src1[30]~q ),
	.datad(!\E_src1[29]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[0]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[0]~18 .extended_lut = "off";
defparam \E_rot_step1[0]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[0]~18 .shared_arith = "off";

dffeas \M_rot_prestep2[4] (
	.clk(clk_clk),
	.d(\E_rot_step1[0]~18_combout ),
	.asdata(\E_rot_step1[4]~19_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[4]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[4] .is_wysiwyg = "true";
defparam \M_rot_prestep2[4] .power_up = "low";

dffeas \M_rot_prestep2[28] (
	.clk(clk_clk),
	.d(\E_rot_step1[24]~20_combout ),
	.asdata(\E_rot_step1[28]~21_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[28]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[28] .is_wysiwyg = "true";
defparam \M_rot_prestep2[28] .power_up = "low";

cyclonev_lcell_comb \M_rot[4]~15 (
	.dataa(!\M_rot_prestep2[20]~q ),
	.datab(!\M_rot_prestep2[12]~q ),
	.datac(!\M_rot_prestep2[4]~q ),
	.datad(!\M_rot_prestep2[28]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~15 .extended_lut = "off";
defparam \M_rot[4]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~15 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~15 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[4]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[4]~15_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~15 .extended_lut = "off";
defparam \A_shift_rot_result~15 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~15 .shared_arith = "off";

dffeas \A_shift_rot_result[20] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~15_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[20]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[20] .is_wysiwyg = "true";
defparam \A_shift_rot_result[20] .power_up = "low";

dffeas \A_slow_inst_result[20] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[20]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[20]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[20] .is_wysiwyg = "true";
defparam \A_slow_inst_result[20] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[20]~35 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[20]~q ),
	.dataf(!\A_slow_inst_result[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[20]~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[20]~35 .extended_lut = "off";
defparam \A_wr_data_unfiltered[20]~35 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[20]~35 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[20]~36 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[20]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[20]~q ),
	.datae(!\A_wr_data_unfiltered[20]~35_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[20]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[20]~36 .extended_lut = "off";
defparam \A_wr_data_unfiltered[20]~36 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[20]~36 .shared_arith = "off";

dffeas \W_wr_data[20] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[20]~36_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[20]~q ),
	.prn(vcc));
defparam \W_wr_data[20] .is_wysiwyg = "true";
defparam \W_wr_data[20] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[20]~25 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[20] ),
	.datab(!\W_wr_data[20]~q ),
	.datac(!\M_alu_result[20]~q ),
	.datad(!\A_wr_data_unfiltered[20]~36_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[20]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[20]~25 .extended_lut = "off";
defparam \D_src1_reg[20]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[20]~25 .shared_arith = "off";

dffeas \E_src1[20] (
	.clk(clk_clk),
	.d(\D_src1_reg[20]~25_combout ),
	.asdata(\E_alu_result[20]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[20]~q ),
	.prn(vcc));
defparam \E_src1[20] .is_wysiwyg = "true";
defparam \E_src1[20] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~15 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[20]~q ),
	.datae(!\E_src1[20]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~15 .extended_lut = "off";
defparam \E_alu_result~15 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~15 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[20]~70 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~15_combout ),
	.datad(!\Add17~77_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[20]~70_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[20]~70 .extended_lut = "off";
defparam \D_src2_reg[20]~70 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[20]~70 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[20]~31 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[20]~q ),
	.datae(!\A_wr_data_unfiltered[20]~36_combout ),
	.dataf(!\M_alu_result[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[20]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[20]~31 .extended_lut = "off";
defparam \D_src2_reg[20]~31 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[20]~31 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[20]~22 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[10]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[20]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[20]~22 .extended_lut = "off";
defparam \D_src2[20]~22 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \D_src2[20]~22 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[20]~23 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[20]~70_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.datae(!\D_src2_reg[20]~31_combout ),
	.dataf(!\D_src2[20]~22_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[20]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[20]~23 .extended_lut = "off";
defparam \D_src2[20]~23 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[20]~23 .shared_arith = "off";

dffeas \E_src2[20] (
	.clk(clk_clk),
	.d(\D_src2[20]~23_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[20]~q ),
	.prn(vcc));
defparam \E_src2[20] .is_wysiwyg = "true";
defparam \E_src2[20] .power_up = "low";

cyclonev_lcell_comb \Add17~73 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[21]~q ),
	.datae(gnd),
	.dataf(!\E_src1[21]~q ),
	.datag(gnd),
	.cin(\Add17~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~73_sumout ),
	.cout(\Add17~74 ),
	.shareout());
defparam \Add17~73 .extended_lut = "off";
defparam \Add17~73 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~73 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[21] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~14_combout ),
	.datac(!\Add17~73_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[21]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[21] .extended_lut = "off";
defparam \E_alu_result[21] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[21] .shared_arith = "off";

dffeas \M_alu_result[21] (
	.clk(clk_clk),
	.d(\E_alu_result[21]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[21]~q ),
	.prn(vcc));
defparam \M_alu_result[21] .is_wysiwyg = "true";
defparam \M_alu_result[21] .power_up = "low";

dffeas \A_inst_result[21] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[21] ),
	.asdata(\M_alu_result[21]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[21]~q ),
	.prn(vcc));
defparam \A_inst_result[21] .is_wysiwyg = "true";
defparam \A_inst_result[21] .power_up = "low";

cyclonev_lcell_comb \M_rot[5]~14 (
	.dataa(!\M_rot_prestep2[21]~q ),
	.datab(!\M_rot_prestep2[13]~q ),
	.datac(!\M_rot_prestep2[5]~q ),
	.datad(!\M_rot_prestep2[29]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~14 .extended_lut = "off";
defparam \M_rot[5]~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~14 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~14 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[5]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[5]~14_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~14 .extended_lut = "off";
defparam \A_shift_rot_result~14 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~14 .shared_arith = "off";

dffeas \A_shift_rot_result[21] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~14_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[21]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[21] .is_wysiwyg = "true";
defparam \A_shift_rot_result[21] .power_up = "low";

dffeas \A_slow_inst_result[21] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[21]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[21]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[21] .is_wysiwyg = "true";
defparam \A_slow_inst_result[21] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[21]~33 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[21]~q ),
	.dataf(!\A_slow_inst_result[21]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[21]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[21]~33 .extended_lut = "off";
defparam \A_wr_data_unfiltered[21]~33 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[21]~33 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[21]~34 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[21]~q ),
	.datac(!\A_mul_result[21]~q ),
	.datad(!\A_wr_data_unfiltered[29]~32_combout ),
	.datae(!\A_wr_data_unfiltered[21]~33_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[21]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[21]~34 .extended_lut = "off";
defparam \A_wr_data_unfiltered[21]~34 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \A_wr_data_unfiltered[21]~34 .shared_arith = "off";

dffeas \W_wr_data[21] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[21]~34_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[21]~q ),
	.prn(vcc));
defparam \W_wr_data[21] .is_wysiwyg = "true";
defparam \W_wr_data[21] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[21]~22 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[21] ),
	.datab(!\W_wr_data[21]~q ),
	.datac(!\M_alu_result[21]~q ),
	.datad(!\A_wr_data_unfiltered[21]~34_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[21]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[21]~22 .extended_lut = "off";
defparam \D_src1_reg[21]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[21]~22 .shared_arith = "off";

dffeas \E_src1[21] (
	.clk(clk_clk),
	.d(\D_src1_reg[21]~22_combout ),
	.asdata(\E_alu_result[21]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[21]~q ),
	.prn(vcc));
defparam \E_src1[21] .is_wysiwyg = "true";
defparam \E_src1[21] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[21]~10 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[21]~q ),
	.datad(!\E_src1[21]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[21]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[21]~10 .extended_lut = "off";
defparam \E_logic_result[21]~10 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[21]~10 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~14 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_result[21]~10_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~14 .extended_lut = "off";
defparam \E_alu_result~14 .lut_mask = 64'h7777777777777777;
defparam \E_alu_result~14 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[21]~68 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~14_combout ),
	.datad(!\Add17~73_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[21]~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[21]~68 .extended_lut = "off";
defparam \D_src2_reg[21]~68 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[21]~68 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[21]~29 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[21]~q ),
	.datae(!\A_wr_data_unfiltered[21]~34_combout ),
	.dataf(!\M_alu_result[21]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[21]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[21]~29 .extended_lut = "off";
defparam \D_src2_reg[21]~29 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[21]~29 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[21]~18 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[21]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[21]~18 .extended_lut = "off";
defparam \D_src2[21]~18 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[21]~18 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[21]~19 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[21]~68_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.datae(!\D_src2_reg[21]~29_combout ),
	.dataf(!\D_src2[21]~18_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[21]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[21]~19 .extended_lut = "off";
defparam \D_src2[21]~19 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[21]~19 .shared_arith = "off";

dffeas \E_src2[21] (
	.clk(clk_clk),
	.d(\D_src2[21]~19_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[21]~q ),
	.prn(vcc));
defparam \E_src2[21] .is_wysiwyg = "true";
defparam \E_src2[21] .power_up = "low";

cyclonev_lcell_comb \Add17~121 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[22]~q ),
	.datae(gnd),
	.dataf(!\E_src1[22]~q ),
	.datag(gnd),
	.cin(\Add17~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~121_sumout ),
	.cout(\Add17~122 ),
	.shareout());
defparam \Add17~121 .extended_lut = "off";
defparam \Add17~121 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~121 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[22] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~26_combout ),
	.datac(!\Add17~121_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[22]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[22] .extended_lut = "off";
defparam \E_alu_result[22] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[22] .shared_arith = "off";

dffeas \M_alu_result[22] (
	.clk(clk_clk),
	.d(\E_alu_result[22]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[22]~q ),
	.prn(vcc));
defparam \M_alu_result[22] .is_wysiwyg = "true";
defparam \M_alu_result[22] .power_up = "low";

dffeas \A_inst_result[22] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[22] ),
	.asdata(\M_alu_result[22]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[22]~q ),
	.prn(vcc));
defparam \A_inst_result[22] .is_wysiwyg = "true";
defparam \A_inst_result[22] .power_up = "low";

cyclonev_lcell_comb \M_rot[6]~26 (
	.dataa(!\M_rot_prestep2[22]~q ),
	.datab(!\M_rot_prestep2[14]~q ),
	.datac(!\M_rot_prestep2[6]~q ),
	.datad(!\M_rot_prestep2[30]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~26 .extended_lut = "off";
defparam \M_rot[6]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~26 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~26 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[6]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[6]~26_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~26 .extended_lut = "off";
defparam \A_shift_rot_result~26 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~26 .shared_arith = "off";

dffeas \A_shift_rot_result[22] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~26_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[22]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[22] .is_wysiwyg = "true";
defparam \A_shift_rot_result[22] .power_up = "low";

dffeas \A_slow_inst_result[22] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[22]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[22]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[22] .is_wysiwyg = "true";
defparam \A_slow_inst_result[22] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[22]~56 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[22]~q ),
	.dataf(!\A_slow_inst_result[22]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[22]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[22]~56 .extended_lut = "off";
defparam \A_wr_data_unfiltered[22]~56 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[22]~56 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[22]~57 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[22]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[22]~q ),
	.datae(!\A_wr_data_unfiltered[22]~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[22]~57_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[22]~57 .extended_lut = "off";
defparam \A_wr_data_unfiltered[22]~57 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[22]~57 .shared_arith = "off";

dffeas \W_wr_data[22] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[22]~57_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[22]~q ),
	.prn(vcc));
defparam \W_wr_data[22] .is_wysiwyg = "true";
defparam \W_wr_data[22] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[22]~26 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\W_wr_data[22]~q ),
	.datac(!\M_alu_result[22]~q ),
	.datad(!\A_wr_data_unfiltered[22]~57_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[22]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[22]~26 .extended_lut = "off";
defparam \D_src1_reg[22]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[22]~26 .shared_arith = "off";

dffeas \E_src1[22] (
	.clk(clk_clk),
	.d(\D_src1_reg[22]~26_combout ),
	.asdata(\E_alu_result[22]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[22]~q ),
	.prn(vcc));
defparam \E_src1[22] .is_wysiwyg = "true";
defparam \E_src1[22] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~26 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[22]~q ),
	.datae(!\E_src1[22]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~26 .extended_lut = "off";
defparam \E_alu_result~26 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~26 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[22]~71 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~26_combout ),
	.datad(!\Add17~121_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[22]~71_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[22]~71 .extended_lut = "off";
defparam \D_src2_reg[22]~71 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[22]~71 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[22]~52 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[22]~q ),
	.datae(!\A_wr_data_unfiltered[22]~57_combout ),
	.dataf(!\M_alu_result[22]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[22]~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[22]~52 .extended_lut = "off";
defparam \D_src2_reg[22]~52 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[22]~52 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[22]~24 (
	.dataa(!\D_iw[12]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[22]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[22]~24 .extended_lut = "off";
defparam \D_src2[22]~24 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[22]~24 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[22]~25 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[22]~71_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.datae(!\D_src2_reg[22]~52_combout ),
	.dataf(!\D_src2[22]~24_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[22]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[22]~25 .extended_lut = "off";
defparam \D_src2[22]~25 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[22]~25 .shared_arith = "off";

dffeas \E_src2[22] (
	.clk(clk_clk),
	.d(\D_src2[22]~25_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[22]~q ),
	.prn(vcc));
defparam \E_src2[22] .is_wysiwyg = "true";
defparam \E_src2[22] .power_up = "low";

cyclonev_lcell_comb \Add17~113 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[23]~q ),
	.datae(gnd),
	.dataf(!\E_src1[23]~q ),
	.datag(gnd),
	.cin(\Add17~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~113_sumout ),
	.cout(\Add17~114 ),
	.shareout());
defparam \Add17~113 .extended_lut = "off";
defparam \Add17~113 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~113 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[23] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~24_combout ),
	.datac(!\Add17~113_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[23]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[23] .extended_lut = "off";
defparam \E_alu_result[23] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[23] .shared_arith = "off";

dffeas \M_alu_result[23] (
	.clk(clk_clk),
	.d(\E_alu_result[23]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[23]~q ),
	.prn(vcc));
defparam \M_alu_result[23] .is_wysiwyg = "true";
defparam \M_alu_result[23] .power_up = "low";

dffeas \A_inst_result[23] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.asdata(\M_alu_result[23]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[23]~q ),
	.prn(vcc));
defparam \A_inst_result[23] .is_wysiwyg = "true";
defparam \A_inst_result[23] .power_up = "low";

cyclonev_lcell_comb \M_rot[7]~24 (
	.dataa(!\M_rot_prestep2[23]~q ),
	.datab(!\M_rot_prestep2[15]~q ),
	.datac(!\M_rot_prestep2[7]~q ),
	.datad(!\M_rot_prestep2[31]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~24 .extended_lut = "off";
defparam \M_rot[7]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~24 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~24 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[7]~q ),
	.datac(!\M_rot_pass2~q ),
	.datad(!\M_rot_sel_fill2~q ),
	.datae(!\M_rot[7]~24_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~24 .extended_lut = "off";
defparam \A_shift_rot_result~24 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~24 .shared_arith = "off";

dffeas \A_shift_rot_result[23] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~24_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[23]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[23] .is_wysiwyg = "true";
defparam \A_shift_rot_result[23] .power_up = "low";

dffeas \A_slow_inst_result[23] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[23]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[23]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[23] .is_wysiwyg = "true";
defparam \A_slow_inst_result[23] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[23]~53 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[23]~q ),
	.dataf(!\A_slow_inst_result[23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[23]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[23]~53 .extended_lut = "off";
defparam \A_wr_data_unfiltered[23]~53 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[23]~53 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[23]~54 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[23]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[23]~q ),
	.datae(!\A_wr_data_unfiltered[23]~53_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[23]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[23]~54 .extended_lut = "off";
defparam \A_wr_data_unfiltered[23]~54 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[23]~54 .shared_arith = "off";

dffeas \W_wr_data[23] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[23]~54_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[23]~q ),
	.prn(vcc));
defparam \W_wr_data[23] .is_wysiwyg = "true";
defparam \W_wr_data[23] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[23]~29 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[23] ),
	.datab(!\W_wr_data[23]~q ),
	.datac(!\M_alu_result[23]~q ),
	.datad(!\A_wr_data_unfiltered[23]~54_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[23]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[23]~29 .extended_lut = "off";
defparam \D_src1_reg[23]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[23]~29 .shared_arith = "off";

dffeas \E_src1[23] (
	.clk(clk_clk),
	.d(\D_src1_reg[23]~29_combout ),
	.asdata(\E_alu_result[23]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[23]~q ),
	.prn(vcc));
defparam \E_src1[23] .is_wysiwyg = "true";
defparam \E_src1[23] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~24 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[23]~q ),
	.datae(!\E_src1[23]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~24 .extended_lut = "off";
defparam \E_alu_result~24 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~24 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[23]~73 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~24_combout ),
	.datad(!\Add17~113_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~73_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~73 .extended_lut = "off";
defparam \D_src2_reg[23]~73 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[23]~73 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[23]~49 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[23]~q ),
	.datae(!\A_wr_data_unfiltered[23]~54_combout ),
	.dataf(!\M_alu_result[23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~49 .extended_lut = "off";
defparam \D_src2_reg[23]~49 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[23]~49 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[23]~28 (
	.dataa(!\D_iw[13]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[23]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[23]~28 .extended_lut = "off";
defparam \D_src2[23]~28 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[23]~28 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[23]~29 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[23]~73_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.datae(!\D_src2_reg[23]~49_combout ),
	.dataf(!\D_src2[23]~28_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[23]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[23]~29 .extended_lut = "off";
defparam \D_src2[23]~29 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[23]~29 .shared_arith = "off";

dffeas \E_src2[23] (
	.clk(clk_clk),
	.d(\D_src2[23]~29_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[23]~q ),
	.prn(vcc));
defparam \E_src2[23] .is_wysiwyg = "true";
defparam \E_src2[23] .power_up = "low";

cyclonev_lcell_comb \Add17~89 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[24]~q ),
	.datae(gnd),
	.dataf(!\E_src1[24]~q ),
	.datag(gnd),
	.cin(\Add17~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~89_sumout ),
	.cout(\Add17~90 ),
	.shareout());
defparam \Add17~89 .extended_lut = "off";
defparam \Add17~89 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~89 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[24] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~18_combout ),
	.datac(!\Add17~89_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[24]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[24] .extended_lut = "off";
defparam \E_alu_result[24] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[24] .shared_arith = "off";

dffeas \M_alu_result[24] (
	.clk(clk_clk),
	.d(\E_alu_result[24]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[24]~q ),
	.prn(vcc));
defparam \M_alu_result[24] .is_wysiwyg = "true";
defparam \M_alu_result[24] .power_up = "low";

dffeas \A_inst_result[24] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[24] ),
	.asdata(\M_alu_result[24]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[24]~q ),
	.prn(vcc));
defparam \A_inst_result[24] .is_wysiwyg = "true";
defparam \A_inst_result[24] .power_up = "low";

cyclonev_lcell_comb \M_rot[0]~18 (
	.dataa(!\M_rot_prestep2[24]~q ),
	.datab(!\M_rot_prestep2[16]~q ),
	.datac(!\M_rot_prestep2[8]~q ),
	.datad(!\M_rot_prestep2[0]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~18 .extended_lut = "off";
defparam \M_rot[0]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~18 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~18 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[0]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[0]~18_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~18 .extended_lut = "off";
defparam \A_shift_rot_result~18 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~18 .shared_arith = "off";

dffeas \A_shift_rot_result[24] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~18_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[24]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[24] .is_wysiwyg = "true";
defparam \A_shift_rot_result[24] .power_up = "low";

dffeas \A_slow_inst_result[24] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[24]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[24]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[24] .is_wysiwyg = "true";
defparam \A_slow_inst_result[24] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[24]~41 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[24]~q ),
	.dataf(!\A_slow_inst_result[24]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[24]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[24]~41 .extended_lut = "off";
defparam \A_wr_data_unfiltered[24]~41 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[24]~41 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[24]~42 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[24]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[24]~q ),
	.datae(!\A_wr_data_unfiltered[24]~41_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[24]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[24]~42 .extended_lut = "off";
defparam \A_wr_data_unfiltered[24]~42 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[24]~42 .shared_arith = "off";

dffeas \W_wr_data[24] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[24]~42_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[24]~q ),
	.prn(vcc));
defparam \W_wr_data[24] .is_wysiwyg = "true";
defparam \W_wr_data[24] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[24]~28 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[24] ),
	.datab(!\W_wr_data[24]~q ),
	.datac(!\M_alu_result[24]~q ),
	.datad(!\A_wr_data_unfiltered[24]~42_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[24]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[24]~28 .extended_lut = "off";
defparam \D_src1_reg[24]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[24]~28 .shared_arith = "off";

dffeas \E_src1[24] (
	.clk(clk_clk),
	.d(\D_src1_reg[24]~28_combout ),
	.asdata(\E_alu_result[24]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[24]~q ),
	.prn(vcc));
defparam \E_src1[24] .is_wysiwyg = "true";
defparam \E_src1[24] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~18 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[24]~q ),
	.datae(!\E_src1[24]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~18 .extended_lut = "off";
defparam \E_alu_result~18 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~18 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[24]~72 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~18_combout ),
	.datad(!\Add17~89_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~72_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~72 .extended_lut = "off";
defparam \D_src2_reg[24]~72 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[24]~72 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[24]~37 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[24]~q ),
	.datae(!\A_wr_data_unfiltered[24]~42_combout ),
	.dataf(!\M_alu_result[24]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~37 .extended_lut = "off";
defparam \D_src2_reg[24]~37 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[24]~37 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[24]~26 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[24]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[24]~26 .extended_lut = "off";
defparam \D_src2[24]~26 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[24]~26 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[24]~27 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[24]~72_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.datae(!\D_src2_reg[24]~37_combout ),
	.dataf(!\D_src2[24]~26_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[24]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[24]~27 .extended_lut = "off";
defparam \D_src2[24]~27 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[24]~27 .shared_arith = "off";

dffeas \E_src2[24] (
	.clk(clk_clk),
	.d(\D_src2[24]~27_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[24]~q ),
	.prn(vcc));
defparam \E_src2[24] .is_wysiwyg = "true";
defparam \E_src2[24] .power_up = "low";

cyclonev_lcell_comb \Add17~81 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[25]~q ),
	.datae(gnd),
	.dataf(!\E_src1[25]~q ),
	.datag(gnd),
	.cin(\Add17~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~81_sumout ),
	.cout(\Add17~82 ),
	.shareout());
defparam \Add17~81 .extended_lut = "off";
defparam \Add17~81 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~81 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[25] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~16_combout ),
	.datac(!\Add17~81_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[25]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[25] .extended_lut = "off";
defparam \E_alu_result[25] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[25] .shared_arith = "off";

dffeas \M_alu_result[25] (
	.clk(clk_clk),
	.d(\E_alu_result[25]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[25]~q ),
	.prn(vcc));
defparam \M_alu_result[25] .is_wysiwyg = "true";
defparam \M_alu_result[25] .power_up = "low";

dffeas \A_inst_result[25] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[25] ),
	.asdata(\M_alu_result[25]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[25]~q ),
	.prn(vcc));
defparam \A_inst_result[25] .is_wysiwyg = "true";
defparam \A_inst_result[25] .power_up = "low";

cyclonev_lcell_comb \M_rot[1]~16 (
	.dataa(!\M_rot_prestep2[25]~q ),
	.datab(!\M_rot_prestep2[17]~q ),
	.datac(!\M_rot_prestep2[9]~q ),
	.datad(!\M_rot_prestep2[1]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~16 .extended_lut = "off";
defparam \M_rot[1]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~16 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~16 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[1]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[1]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~16 .extended_lut = "off";
defparam \A_shift_rot_result~16 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~16 .shared_arith = "off";

dffeas \A_shift_rot_result[25] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~16_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[25]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[25] .is_wysiwyg = "true";
defparam \A_shift_rot_result[25] .power_up = "low";

dffeas \A_slow_inst_result[25] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[25]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[25]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[25] .is_wysiwyg = "true";
defparam \A_slow_inst_result[25] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[25]~37 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[25]~q ),
	.dataf(!\A_slow_inst_result[25]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[25]~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[25]~37 .extended_lut = "off";
defparam \A_wr_data_unfiltered[25]~37 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[25]~37 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[25]~38 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[25]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[25]~q ),
	.datae(!\A_wr_data_unfiltered[25]~37_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[25]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[25]~38 .extended_lut = "off";
defparam \A_wr_data_unfiltered[25]~38 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[25]~38 .shared_arith = "off";

dffeas \W_wr_data[25] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[25]~38_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[25]~q ),
	.prn(vcc));
defparam \W_wr_data[25] .is_wysiwyg = "true";
defparam \W_wr_data[25] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[25]~24 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[25] ),
	.datab(!\W_wr_data[25]~q ),
	.datac(!\M_alu_result[25]~q ),
	.datad(!\A_wr_data_unfiltered[25]~38_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[25]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[25]~24 .extended_lut = "off";
defparam \D_src1_reg[25]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[25]~24 .shared_arith = "off";

dffeas \E_src1[25] (
	.clk(clk_clk),
	.d(\D_src1_reg[25]~24_combout ),
	.asdata(\E_alu_result[25]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[25]~q ),
	.prn(vcc));
defparam \E_src1[25] .is_wysiwyg = "true";
defparam \E_src1[25] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~16 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[25]~q ),
	.datae(!\E_src1[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~16 .extended_lut = "off";
defparam \E_alu_result~16 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~16 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[25]~69 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~16_combout ),
	.datad(!\Add17~81_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~69_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~69 .extended_lut = "off";
defparam \D_src2_reg[25]~69 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[25]~69 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[25]~33 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[25]~q ),
	.datae(!\A_wr_data_unfiltered[25]~38_combout ),
	.dataf(!\M_alu_result[25]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~33 .extended_lut = "off";
defparam \D_src2_reg[25]~33 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[25]~33 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[25]~20 (
	.dataa(!\D_iw[15]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[25]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[25]~20 .extended_lut = "off";
defparam \D_src2[25]~20 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[25]~20 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[25]~21 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[25]~69_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.datae(!\D_src2_reg[25]~33_combout ),
	.dataf(!\D_src2[25]~20_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[25]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[25]~21 .extended_lut = "off";
defparam \D_src2[25]~21 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[25]~21 .shared_arith = "off";

dffeas \E_src2[25] (
	.clk(clk_clk),
	.d(\D_src2[25]~21_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[25]~q ),
	.prn(vcc));
defparam \E_src2[25] .is_wysiwyg = "true";
defparam \E_src2[25] .power_up = "low";

cyclonev_lcell_comb \Add17~105 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[26]~q ),
	.datae(gnd),
	.dataf(!\E_src1[26]~q ),
	.datag(gnd),
	.cin(\Add17~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~105_sumout ),
	.cout(\Add17~106 ),
	.shareout());
defparam \Add17~105 .extended_lut = "off";
defparam \Add17~105 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~105 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[26] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~22_combout ),
	.datac(!\Add17~105_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[26]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[26] .extended_lut = "off";
defparam \E_alu_result[26] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[26] .shared_arith = "off";

dffeas \M_alu_result[26] (
	.clk(clk_clk),
	.d(\E_alu_result[26]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[26]~q ),
	.prn(vcc));
defparam \M_alu_result[26] .is_wysiwyg = "true";
defparam \M_alu_result[26] .power_up = "low";

dffeas \A_inst_result[26] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[26] ),
	.asdata(\M_alu_result[26]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[26]~q ),
	.prn(vcc));
defparam \A_inst_result[26] .is_wysiwyg = "true";
defparam \A_inst_result[26] .power_up = "low";

cyclonev_lcell_comb \M_rot[2]~22 (
	.dataa(!\M_rot_prestep2[26]~q ),
	.datab(!\M_rot_prestep2[18]~q ),
	.datac(!\M_rot_prestep2[10]~q ),
	.datad(!\M_rot_prestep2[2]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~22 .extended_lut = "off";
defparam \M_rot[2]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~22 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~22 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[2]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[2]~22_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~22 .extended_lut = "off";
defparam \A_shift_rot_result~22 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~22 .shared_arith = "off";

dffeas \A_shift_rot_result[26] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~22_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[26]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[26] .is_wysiwyg = "true";
defparam \A_shift_rot_result[26] .power_up = "low";

dffeas \A_slow_inst_result[26] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[26]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[26]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[26] .is_wysiwyg = "true";
defparam \A_slow_inst_result[26] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[26]~49 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[26]~q ),
	.dataf(!\A_slow_inst_result[26]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[26]~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[26]~49 .extended_lut = "off";
defparam \A_wr_data_unfiltered[26]~49 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[26]~49 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[26]~50 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[26]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[26]~q ),
	.datae(!\A_wr_data_unfiltered[26]~49_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[26]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[26]~50 .extended_lut = "off";
defparam \A_wr_data_unfiltered[26]~50 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[26]~50 .shared_arith = "off";

dffeas \W_wr_data[26] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[26]~50_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[26]~q ),
	.prn(vcc));
defparam \W_wr_data[26] .is_wysiwyg = "true";
defparam \W_wr_data[26] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[26]~20 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[26] ),
	.datab(!\W_wr_data[26]~q ),
	.datac(!\M_alu_result[26]~q ),
	.datad(!\A_wr_data_unfiltered[26]~50_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[26]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[26]~20 .extended_lut = "off";
defparam \D_src1_reg[26]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[26]~20 .shared_arith = "off";

dffeas \E_src1[26] (
	.clk(clk_clk),
	.d(\D_src1_reg[26]~20_combout ),
	.asdata(\E_alu_result[26]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[26]~q ),
	.prn(vcc));
defparam \E_src1[26] .is_wysiwyg = "true";
defparam \E_src1[26] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~22 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[26]~q ),
	.datae(!\E_src1[26]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~22 .extended_lut = "off";
defparam \E_alu_result~22 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~22 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[26]~66 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~22_combout ),
	.datad(!\Add17~105_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~66 .extended_lut = "off";
defparam \D_src2_reg[26]~66 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[26]~66 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[26]~45 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[26]~q ),
	.datae(!\A_wr_data_unfiltered[26]~50_combout ),
	.dataf(!\M_alu_result[26]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~45 .extended_lut = "off";
defparam \D_src2_reg[26]~45 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[26]~45 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[26]~14 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_ctrl_hi_imm16~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[26]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[26]~14 .extended_lut = "off";
defparam \D_src2[26]~14 .lut_mask = 64'h7FDF7FDF7FDF7FDF;
defparam \D_src2[26]~14 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[26]~15 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[26]~66_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.datae(!\D_src2_reg[26]~45_combout ),
	.dataf(!\D_src2[26]~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[26]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[26]~15 .extended_lut = "off";
defparam \D_src2[26]~15 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[26]~15 .shared_arith = "off";

dffeas \E_src2[26] (
	.clk(clk_clk),
	.d(\D_src2[26]~15_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[26]~q ),
	.prn(vcc));
defparam \E_src2[26] .is_wysiwyg = "true";
defparam \E_src2[26] .power_up = "low";

cyclonev_lcell_comb \Add17~97 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[27]~q ),
	.datae(gnd),
	.dataf(!\E_src1[27]~q ),
	.datag(gnd),
	.cin(\Add17~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~97_sumout ),
	.cout(\Add17~98 ),
	.shareout());
defparam \Add17~97 .extended_lut = "off";
defparam \Add17~97 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~97 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[28]~63 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~31_combout ),
	.datad(!\Add17~133_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~63 .extended_lut = "off";
defparam \D_src2_reg[28]~63 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[28]~63 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[28]~64 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[28]~q ),
	.datae(!\A_wr_data_unfiltered[28]~66_combout ),
	.dataf(!\M_alu_result[28]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~64 .extended_lut = "off";
defparam \D_src2_reg[28]~64 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[28]~64 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[28]~10 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[18]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[28]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[28]~10 .extended_lut = "off";
defparam \D_src2[28]~10 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \D_src2[28]~10 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[28]~11 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[28]~63_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.datae(!\D_src2_reg[28]~64_combout ),
	.dataf(!\D_src2[28]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[28]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[28]~11 .extended_lut = "off";
defparam \D_src2[28]~11 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[28]~11 .shared_arith = "off";

dffeas \E_src2[28] (
	.clk(clk_clk),
	.d(\D_src2[28]~11_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[28]~q ),
	.prn(vcc));
defparam \E_src2[28] .is_wysiwyg = "true";
defparam \E_src2[28] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~31 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[28]~q ),
	.datae(!\E_src1[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~31 .extended_lut = "off";
defparam \E_alu_result~31 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~31 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[28] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~31_combout ),
	.datac(!\Add17~133_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[28]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[28] .extended_lut = "off";
defparam \E_alu_result[28] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[28] .shared_arith = "off";

dffeas \M_alu_result[28] (
	.clk(clk_clk),
	.d(\E_alu_result[28]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[28]~q ),
	.prn(vcc));
defparam \M_alu_result[28] .is_wysiwyg = "true";
defparam \M_alu_result[28] .power_up = "low";

dffeas \A_inst_result[28] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[28] ),
	.asdata(\M_alu_result[28]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[28]~q ),
	.prn(vcc));
defparam \A_inst_result[28] .is_wysiwyg = "true";
defparam \A_inst_result[28] .power_up = "low";

cyclonev_lcell_comb \M_rot[4]~31 (
	.dataa(!\M_rot_prestep2[28]~q ),
	.datab(!\M_rot_prestep2[20]~q ),
	.datac(!\M_rot_prestep2[12]~q ),
	.datad(!\M_rot_prestep2[4]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~31 .extended_lut = "off";
defparam \M_rot[4]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~31 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~31 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[4]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[4]~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~31 .extended_lut = "off";
defparam \A_shift_rot_result~31 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~31 .shared_arith = "off";

dffeas \A_shift_rot_result[28] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~31_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[28]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[28] .is_wysiwyg = "true";
defparam \A_shift_rot_result[28] .power_up = "low";

dffeas \A_slow_inst_result[28] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[28]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[28]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[28] .is_wysiwyg = "true";
defparam \A_slow_inst_result[28] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[28]~65 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[28]~q ),
	.dataf(!\A_slow_inst_result[28]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[28]~65_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[28]~65 .extended_lut = "off";
defparam \A_wr_data_unfiltered[28]~65 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[28]~65 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[28]~66 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[28]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[28]~q ),
	.datae(!\A_wr_data_unfiltered[28]~65_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[28]~66_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[28]~66 .extended_lut = "off";
defparam \A_wr_data_unfiltered[28]~66 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[28]~66 .shared_arith = "off";

dffeas \W_wr_data[28] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[28]~66_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[28]~q ),
	.prn(vcc));
defparam \W_wr_data[28] .is_wysiwyg = "true";
defparam \W_wr_data[28] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[28]~18 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[28] ),
	.datab(!\W_wr_data[28]~q ),
	.datac(!\M_alu_result[28]~q ),
	.datad(!\A_wr_data_unfiltered[28]~66_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[28]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[28]~18 .extended_lut = "off";
defparam \D_src1_reg[28]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[28]~18 .shared_arith = "off";

dffeas \E_src1[28] (
	.clk(clk_clk),
	.d(\D_src1_reg[28]~18_combout ),
	.asdata(\E_alu_result[28]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[28]~q ),
	.prn(vcc));
defparam \E_src1[28] .is_wysiwyg = "true";
defparam \E_src1[28] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[28]~21 (
	.dataa(!\E_src1[28]~q ),
	.datab(!\E_src1[27]~q ),
	.datac(!\E_src1[26]~q ),
	.datad(!\E_src1[25]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[28]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[28]~21 .extended_lut = "off";
defparam \E_rot_step1[28]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[28]~21 .shared_arith = "off";

dffeas \M_rot_prestep2[0] (
	.clk(clk_clk),
	.d(\E_rot_step1[28]~21_combout ),
	.asdata(\E_rot_step1[0]~18_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[0]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[0] .is_wysiwyg = "true";
defparam \M_rot_prestep2[0] .power_up = "low";

cyclonev_lcell_comb \M_rot[0]~6 (
	.dataa(!\M_rot_prestep2[8]~q ),
	.datab(!\M_rot_prestep2[0]~q ),
	.datac(!\M_rot_prestep2[24]~q ),
	.datad(!\M_rot_prestep2[16]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~6 .extended_lut = "off";
defparam \M_rot[0]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~6 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~6 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_sel_fill1~q ),
	.datad(!\M_rot_mask[0]~q ),
	.datae(!\M_rot[0]~6_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~6 .extended_lut = "off";
defparam \A_shift_rot_result~6 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~6 .shared_arith = "off";

dffeas \A_shift_rot_result[8] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[8]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[8] .is_wysiwyg = "true";
defparam \A_shift_rot_result[8] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte1_data_aligned_nxt[0]~5 (
	.dataa(!\A_ld_align_sh16~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!\d_readdata_d1[24]~q ),
	.datae(!\d_readdata_d1[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte1_data_aligned_nxt[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte1_data_aligned_nxt[0]~5 .extended_lut = "off";
defparam \A_slow_ld_byte1_data_aligned_nxt[0]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_slow_ld_byte1_data_aligned_nxt[0]~5 .shared_arith = "off";

dffeas \A_slow_inst_result[8] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte1_data_aligned_nxt[0]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[8]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[8] .is_wysiwyg = "true";
defparam \A_slow_inst_result[8] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[8]~16 (
	.dataa(!\A_inst_result[8]~q ),
	.datab(!\A_inst_result[24]~q ),
	.datac(!\A_slow_inst_result[8]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[11]~4_combout ),
	.dataf(!\A_wr_data_unfiltered[11]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[8]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[8]~16 .extended_lut = "off";
defparam \A_wr_data_unfiltered[8]~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[8]~16 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[8]~17 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[8]~q ),
	.datad(!\A_shift_rot_result[8]~q ),
	.datae(!\A_wr_data_unfiltered[8]~16_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[8]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[8]~17 .extended_lut = "off";
defparam \A_wr_data_unfiltered[8]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[8]~17 .shared_arith = "off";

dffeas \W_wr_data[8] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[8]~17_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[8]~q ),
	.prn(vcc));
defparam \W_wr_data[8] .is_wysiwyg = "true";
defparam \W_wr_data[8] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[8]~13 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\A_mul_result[8]~q ),
	.datae(!\A_shift_rot_result[8]~q ),
	.dataf(!\A_wr_data_unfiltered[8]~16_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[8]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[8]~13 .extended_lut = "off";
defparam \D_src2_reg[8]~13 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[8]~13 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[8]~97 (
	.dataa(!\M_alu_result[8]~q ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[5]~3_combout ),
	.datad(!\D_src2_reg[13]~8_combout ),
	.datae(!\W_wr_data[8]~q ),
	.dataf(!\D_src2_reg[8]~13_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[8]~97_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[8]~97 .extended_lut = "off";
defparam \D_src2_reg[8]~97 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[8]~97 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[8]~5 (
	.dataa(!\E_src2[8]~q ),
	.datab(!\E_src1[8]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[8]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[8]~5 .extended_lut = "off";
defparam \E_logic_result[8]~5 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[8]~5 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[8]~7 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[8]~5_combout ),
	.datad(!\E_extra_pc[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[8]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[8]~7 .extended_lut = "off";
defparam \E_alu_result[8]~7 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[8]~7 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[8]~108 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[8] ),
	.datad(!\D_src2_reg[8]~97_combout ),
	.datae(!\D_src2_reg[5]~2_combout ),
	.dataf(!\E_alu_result[8]~7_combout ),
	.datag(!\Add17~1_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[8]~108_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[8]~108 .extended_lut = "on";
defparam \D_src2_reg[8]~108 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[8]~108 .shared_arith = "off";

dffeas \E_src2[8] (
	.clk(clk_clk),
	.d(\D_iw[14]~q ),
	.asdata(\D_src2_reg[8]~108_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[8]~q ),
	.prn(vcc));
defparam \E_src2[8] .is_wysiwyg = "true";
defparam \E_src2[8] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[8] (
	.dataa(!\Add17~1_sumout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\E_alu_result[8]~7_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[8]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[8] .extended_lut = "off";
defparam \E_alu_result[8] .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \E_alu_result[8] .shared_arith = "off";

dffeas \M_alu_result[8] (
	.clk(clk_clk),
	.d(\E_alu_result[8]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[8]~q ),
	.prn(vcc));
defparam \M_alu_result[8] .is_wysiwyg = "true";
defparam \M_alu_result[8] .power_up = "low";

dffeas \A_inst_result[8] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[8] ),
	.asdata(\M_alu_result[8]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[8]~q ),
	.prn(vcc));
defparam \A_inst_result[8] .is_wysiwyg = "true";
defparam \A_inst_result[8] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[0]~30 (
	.dataa(!\A_inst_result[0]~q ),
	.datab(!\A_inst_result[8]~q ),
	.datac(!\A_inst_result[16]~q ),
	.datad(!\A_inst_result[24]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[0]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[0]~30 .extended_lut = "off";
defparam \A_wr_data_unfiltered[0]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[0]~30 .shared_arith = "off";

cyclonev_lcell_comb \E_rot_pass0~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass0~0 .extended_lut = "off";
defparam \E_rot_pass0~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \E_rot_pass0~0 .shared_arith = "off";

dffeas M_rot_pass0(
	.clk(clk_clk),
	.d(\E_rot_pass0~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_pass0~q ),
	.prn(vcc));
defparam M_rot_pass0.is_wysiwyg = "true";
defparam M_rot_pass0.power_up = "low";

cyclonev_lcell_comb \E_rot_sel_fill0~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_shift_rot_left~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_sel_fill0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_sel_fill0~0 .extended_lut = "off";
defparam \E_rot_sel_fill0~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_rot_sel_fill0~0 .shared_arith = "off";

dffeas M_rot_sel_fill0(
	.clk(clk_clk),
	.d(\E_rot_sel_fill0~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_sel_fill0~q ),
	.prn(vcc));
defparam M_rot_sel_fill0.is_wysiwyg = "true";
defparam M_rot_sel_fill0.power_up = "low";

cyclonev_lcell_comb \M_rot[0]~13 (
	.dataa(!\M_rot_prestep2[0]~q ),
	.datab(!\M_rot_prestep2[24]~q ),
	.datac(!\M_rot_prestep2[16]~q ),
	.datad(!\M_rot_prestep2[8]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[0]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[0]~13 .extended_lut = "off";
defparam \M_rot[0]~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[0]~13 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~13 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[0]~q ),
	.datac(!\M_rot_pass0~q ),
	.datad(!\M_rot_sel_fill0~q ),
	.datae(!\M_rot[0]~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~13 .extended_lut = "off";
defparam \A_shift_rot_result~13 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~13 .shared_arith = "off";

dffeas \A_shift_rot_result[0] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~13_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[0]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[0] .is_wysiwyg = "true";
defparam \A_shift_rot_result[0] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[0]~1 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_slow_inst_sel~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[0]~1 .extended_lut = "off";
defparam \A_wr_data_unfiltered[0]~1 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \A_wr_data_unfiltered[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[0]~2 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[0]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[0]~2 .extended_lut = "off";
defparam \A_wr_data_unfiltered[0]~2 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_wr_data_unfiltered[0]~2 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[0]~31 (
	.dataa(!\A_slow_inst_result[0]~q ),
	.datab(!\A_wr_data_unfiltered[0]~30_combout ),
	.datac(!\A_mul_result[0]~q ),
	.datad(!\A_shift_rot_result[0]~q ),
	.datae(!\A_wr_data_unfiltered[0]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[0]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[0]~31 .extended_lut = "off";
defparam \A_wr_data_unfiltered[0]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[0]~31 .shared_arith = "off";

dffeas \W_wr_data[0] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[0]~31_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[0]~q ),
	.prn(vcc));
defparam \W_wr_data[0] .is_wysiwyg = "true";
defparam \W_wr_data[0] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[0]~31 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[0] ),
	.datab(!\W_wr_data[0]~q ),
	.datac(!\M_alu_result[0]~q ),
	.datad(!\A_wr_data_unfiltered[0]~31_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[0]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[0]~31 .extended_lut = "off";
defparam \D_src1_reg[0]~31 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[0]~31 .shared_arith = "off";

dffeas \E_src1[0] (
	.clk(clk_clk),
	.d(\D_src1_reg[0]~31_combout ),
	.asdata(\E_alu_result[0]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[0]~q ),
	.prn(vcc));
defparam \E_src1[0] .is_wysiwyg = "true";
defparam \E_src1[0] .power_up = "low";

cyclonev_lcell_comb \Add17~70 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add17~70_cout ),
	.shareout());
defparam \Add17~70 .extended_lut = "off";
defparam \Add17~70 .lut_mask = 64'h0000000000005555;
defparam \Add17~70 .shared_arith = "off";

cyclonev_lcell_comb \Add17~57 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[0]~q ),
	.datae(gnd),
	.dataf(!\E_src1[0]~q ),
	.datag(gnd),
	.cin(\Add17~70_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~57_sumout ),
	.cout(\Add17~58 ),
	.shareout());
defparam \Add17~57 .extended_lut = "off";
defparam \Add17~57 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~57 .shared_arith = "off";

cyclonev_lcell_comb \Add17~53 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[1]~q ),
	.datae(gnd),
	.dataf(!\E_src1[1]~q ),
	.datag(gnd),
	.cin(\Add17~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~53_sumout ),
	.cout(\Add17~54 ),
	.shareout());
defparam \Add17~53 .extended_lut = "off";
defparam \Add17~53 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~53 .shared_arith = "off";

cyclonev_lcell_comb \Add17~25 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[2]~q ),
	.datae(gnd),
	.dataf(!\E_src1[2]~q ),
	.datag(gnd),
	.cin(\Add17~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~25_sumout ),
	.cout(\Add17~26 ),
	.shareout());
defparam \Add17~25 .extended_lut = "off";
defparam \Add17~25 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~25 .shared_arith = "off";

cyclonev_lcell_comb \Add17~29 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[3]~q ),
	.datae(gnd),
	.dataf(!\E_src1[3]~q ),
	.datag(gnd),
	.cin(\Add17~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~29_sumout ),
	.cout(\Add17~30 ),
	.shareout());
defparam \Add17~29 .extended_lut = "off";
defparam \Add17~29 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~29 .shared_arith = "off";

cyclonev_lcell_comb \Add17~33 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[4]~q ),
	.datae(gnd),
	.dataf(!\E_src1[4]~q ),
	.datag(gnd),
	.cin(\Add17~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~33_sumout ),
	.cout(\Add17~34 ),
	.shareout());
defparam \Add17~33 .extended_lut = "off";
defparam \Add17~33 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~33 .shared_arith = "off";

cyclonev_lcell_comb \Add17~17 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[5]~q ),
	.datae(gnd),
	.dataf(!\E_src1[5]~q ),
	.datag(gnd),
	.cin(\Add17~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~17_sumout ),
	.cout(\Add17~18 ),
	.shareout());
defparam \Add17~17 .extended_lut = "off";
defparam \Add17~17 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~17 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~10 (
	.dataa(!\E_src2[5]~q ),
	.datab(!\E_src1[5]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~10 .extended_lut = "off";
defparam \E_alu_result~10 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~10 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[5] (
	.dataa(!\Add17~17_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~10_combout ),
	.datae(!\E_extra_pc[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[5]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[5] .extended_lut = "off";
defparam \E_alu_result[5] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[5] .shared_arith = "off";

dffeas \M_alu_result[5] (
	.clk(clk_clk),
	.d(\E_alu_result[5]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[5]~q ),
	.prn(vcc));
defparam \M_alu_result[5] .is_wysiwyg = "true";
defparam \M_alu_result[5] .power_up = "low";

dffeas \A_inst_result[5] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[5] ),
	.asdata(\M_alu_result[5]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[5]~q ),
	.prn(vcc));
defparam \A_inst_result[5] .is_wysiwyg = "true";
defparam \A_inst_result[5] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[5]~22 (
	.dataa(!\A_inst_result[5]~q ),
	.datab(!\A_inst_result[13]~q ),
	.datac(!\A_inst_result[21]~q ),
	.datad(!\A_inst_result[29]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[5]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[5]~22 .extended_lut = "off";
defparam \A_wr_data_unfiltered[5]~22 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[5]~22 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[5]~9 (
	.dataa(!\M_rot_prestep2[5]~q ),
	.datab(!\M_rot_prestep2[29]~q ),
	.datac(!\M_rot_prestep2[21]~q ),
	.datad(!\M_rot_prestep2[13]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[5]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[5]~9 .extended_lut = "off";
defparam \M_rot[5]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[5]~9 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~9 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[5]~q ),
	.datac(!\M_rot_pass0~q ),
	.datad(!\M_rot_sel_fill0~q ),
	.datae(!\M_rot[5]~9_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~9 .extended_lut = "off";
defparam \A_shift_rot_result~9 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~9 .shared_arith = "off";

dffeas \A_shift_rot_result[5] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~9_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[5]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[5] .is_wysiwyg = "true";
defparam \A_shift_rot_result[5] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[5]~23 (
	.dataa(!\A_slow_inst_result[5]~q ),
	.datab(!\A_wr_data_unfiltered[5]~22_combout ),
	.datac(!\A_mul_result[5]~q ),
	.datad(!\A_shift_rot_result[5]~q ),
	.datae(!\A_wr_data_unfiltered[0]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[5]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[5]~23 .extended_lut = "off";
defparam \A_wr_data_unfiltered[5]~23 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[5]~23 .shared_arith = "off";

dffeas \W_wr_data[5] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[5]~23_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[5]~q ),
	.prn(vcc));
defparam \W_wr_data[5] .is_wysiwyg = "true";
defparam \W_wr_data[5] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[5]~9 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[5] ),
	.datab(!\W_wr_data[5]~q ),
	.datac(!\M_alu_result[5]~q ),
	.datad(!\A_wr_data_unfiltered[5]~23_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[5]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[5]~9 .extended_lut = "off";
defparam \D_src1_reg[5]~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[5]~9 .shared_arith = "off";

dffeas \E_src1[5] (
	.clk(clk_clk),
	.d(\D_src1_reg[5]~9_combout ),
	.asdata(\E_alu_result[5]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[5]~q ),
	.prn(vcc));
defparam \E_src1[5] .is_wysiwyg = "true";
defparam \E_src1[5] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[6]~6 (
	.dataa(!\E_src1[6]~q ),
	.datab(!\E_src1[5]~q ),
	.datac(!\E_src1[4]~q ),
	.datad(!\E_src1[3]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[6]~6 .extended_lut = "off";
defparam \E_rot_step1[6]~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[6]~6 .shared_arith = "off";

dffeas \M_rot_prestep2[10] (
	.clk(clk_clk),
	.d(\E_rot_step1[6]~6_combout ),
	.asdata(\E_rot_step1[10]~7_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[10]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[10] .is_wysiwyg = "true";
defparam \M_rot_prestep2[10] .power_up = "low";

cyclonev_lcell_comb \M_rot[2]~4 (
	.dataa(!\M_rot_prestep2[10]~q ),
	.datab(!\M_rot_prestep2[2]~q ),
	.datac(!\M_rot_prestep2[26]~q ),
	.datad(!\M_rot_prestep2[18]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~4 .extended_lut = "off";
defparam \M_rot[2]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~4 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~4 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_sel_fill1~q ),
	.datad(!\M_rot_mask[2]~q ),
	.datae(!\M_rot[2]~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~4 .extended_lut = "off";
defparam \A_shift_rot_result~4 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~4 .shared_arith = "off";

dffeas \A_shift_rot_result[10] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[10]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[10] .is_wysiwyg = "true";
defparam \A_shift_rot_result[10] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[10]~13 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[10]~q ),
	.datad(!\A_shift_rot_result[10]~q ),
	.datae(!\A_wr_data_unfiltered[10]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[10]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[10]~13 .extended_lut = "off";
defparam \A_wr_data_unfiltered[10]~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[10]~13 .shared_arith = "off";

dffeas \W_wr_data[10] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[10]~13_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[10]~q ),
	.prn(vcc));
defparam \W_wr_data[10] .is_wysiwyg = "true";
defparam \W_wr_data[10] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[10]~4 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[10] ),
	.datab(!\W_wr_data[10]~q ),
	.datac(!\M_alu_result[10]~q ),
	.datad(!\A_wr_data_unfiltered[10]~13_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[10]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[10]~4 .extended_lut = "off";
defparam \D_src1_reg[10]~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[10]~4 .shared_arith = "off";

dffeas \E_src1[10] (
	.clk(clk_clk),
	.d(\D_src1_reg[10]~4_combout ),
	.asdata(\E_alu_result[10]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[10]~q ),
	.prn(vcc));
defparam \E_src1[10] .is_wysiwyg = "true";
defparam \E_src1[10] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[10]~7 (
	.dataa(!\E_src1[10]~q ),
	.datab(!\E_src1[9]~q ),
	.datac(!\E_src1[8]~q ),
	.datad(!\E_src1[7]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[10]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[10]~7 .extended_lut = "off";
defparam \E_rot_step1[10]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[10]~7 .shared_arith = "off";

dffeas \M_rot_prestep2[14] (
	.clk(clk_clk),
	.d(\E_rot_step1[10]~7_combout ),
	.asdata(\E_rot_step1[14]~4_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[14]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[14] .is_wysiwyg = "true";
defparam \M_rot_prestep2[14] .power_up = "low";

cyclonev_lcell_comb \M_rot[6]~27 (
	.dataa(!\M_rot_prestep2[14]~q ),
	.datab(!\M_rot_prestep2[6]~q ),
	.datac(!\M_rot_prestep2[30]~q ),
	.datad(!\M_rot_prestep2[22]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~27 .extended_lut = "off";
defparam \M_rot[6]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~27 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~27 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_sel_fill1~q ),
	.datad(!\M_rot_mask[6]~q ),
	.datae(!\M_rot[6]~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~27 .extended_lut = "off";
defparam \A_shift_rot_result~27 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~27 .shared_arith = "off";

dffeas \A_shift_rot_result[14] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~27_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[14]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[14] .is_wysiwyg = "true";
defparam \A_shift_rot_result[14] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte1_data_aligned_nxt[6]~7 (
	.dataa(!\A_ld_align_sh16~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!\d_readdata_d1[14]~q ),
	.datae(!\d_readdata_d1[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte1_data_aligned_nxt[6]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte1_data_aligned_nxt[6]~7 .extended_lut = "off";
defparam \A_slow_ld_byte1_data_aligned_nxt[6]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_slow_ld_byte1_data_aligned_nxt[6]~7 .shared_arith = "off";

dffeas \A_slow_inst_result[14] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte1_data_aligned_nxt[6]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[14]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[14] .is_wysiwyg = "true";
defparam \A_slow_inst_result[14] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[14]~58 (
	.dataa(!\A_inst_result[14]~q ),
	.datab(!\A_inst_result[30]~q ),
	.datac(!\A_slow_inst_result[14]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[11]~4_combout ),
	.dataf(!\A_wr_data_unfiltered[11]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[14]~58_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[14]~58 .extended_lut = "off";
defparam \A_wr_data_unfiltered[14]~58 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[14]~58 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[14]~68 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[14]~q ),
	.datad(!\A_shift_rot_result[14]~q ),
	.datae(!\A_wr_data_unfiltered[14]~58_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[14]~68_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[14]~68 .extended_lut = "off";
defparam \A_wr_data_unfiltered[14]~68 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[14]~68 .shared_arith = "off";

dffeas \W_wr_data[14] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[14]~68_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[14]~q ),
	.prn(vcc));
defparam \W_wr_data[14] .is_wysiwyg = "true";
defparam \W_wr_data[14] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[14]~54 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\A_mul_result[14]~q ),
	.datae(!\A_shift_rot_result[14]~q ),
	.dataf(!\A_wr_data_unfiltered[14]~58_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[14]~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[14]~54 .extended_lut = "off";
defparam \D_src2_reg[14]~54 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[14]~54 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[14]~99 (
	.dataa(!\D_src2_reg[5]~4_combout ),
	.datab(!\M_alu_result[14]~q ),
	.datac(!\D_src2_reg[5]~3_combout ),
	.datad(!\D_src2_reg[13]~8_combout ),
	.datae(!\W_wr_data[14]~q ),
	.dataf(!\D_src2_reg[14]~54_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[14]~99_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[14]~99 .extended_lut = "off";
defparam \D_src2_reg[14]~99 .lut_mask = 64'hA3FFFFFFFFFFFFFF;
defparam \D_src2_reg[14]~99 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[14]~100 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[14] ),
	.datad(!\D_src2_reg[14]~99_combout ),
	.datae(!\D_src2_reg[5]~2_combout ),
	.dataf(!\Add17~125_sumout ),
	.datag(!\E_alu_result~27_combout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[14]~100_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[14]~100 .extended_lut = "on";
defparam \D_src2_reg[14]~100 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[14]~100 .shared_arith = "off";

dffeas \E_src2[14] (
	.clk(clk_clk),
	.d(\D_iw[20]~q ),
	.asdata(\D_src2_reg[14]~100_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[14]~q ),
	.prn(vcc));
defparam \E_src2[14] .is_wysiwyg = "true";
defparam \E_src2[14] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~27 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_logic_op[1]~q ),
	.datac(!\E_logic_op[0]~q ),
	.datad(!\E_src2[14]~q ),
	.datae(!\E_src1[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~27 .extended_lut = "off";
defparam \E_alu_result~27 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \E_alu_result~27 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[14] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\E_alu_result~27_combout ),
	.datac(!\Add17~125_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[14]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[14] .extended_lut = "off";
defparam \E_alu_result[14] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[14] .shared_arith = "off";

dffeas \M_alu_result[14] (
	.clk(clk_clk),
	.d(\E_alu_result[14]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[14]~q ),
	.prn(vcc));
defparam \M_alu_result[14] .is_wysiwyg = "true";
defparam \M_alu_result[14] .power_up = "low";

dffeas \A_inst_result[14] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[14] ),
	.asdata(\M_alu_result[14]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[14]~q ),
	.prn(vcc));
defparam \A_inst_result[14] .is_wysiwyg = "true";
defparam \A_inst_result[14] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[6]~20 (
	.dataa(!\A_inst_result[6]~q ),
	.datab(!\A_inst_result[14]~q ),
	.datac(!\A_inst_result[22]~q ),
	.datad(!\A_inst_result[30]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[6]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[6]~20 .extended_lut = "off";
defparam \A_wr_data_unfiltered[6]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[6]~20 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[6]~8 (
	.dataa(!\M_rot_prestep2[6]~q ),
	.datab(!\M_rot_prestep2[30]~q ),
	.datac(!\M_rot_prestep2[22]~q ),
	.datad(!\M_rot_prestep2[14]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[6]~8 .extended_lut = "off";
defparam \M_rot[6]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[6]~8 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~8 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_sel_fill0~q ),
	.datad(!\M_rot_mask[6]~q ),
	.datae(!\M_rot[6]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~8 .extended_lut = "off";
defparam \A_shift_rot_result~8 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~8 .shared_arith = "off";

dffeas \A_shift_rot_result[6] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~8_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[6]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[6] .is_wysiwyg = "true";
defparam \A_shift_rot_result[6] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[6]~21 (
	.dataa(!\A_slow_inst_result[6]~q ),
	.datab(!\A_wr_data_unfiltered[6]~20_combout ),
	.datac(!\A_mul_result[6]~q ),
	.datad(!\A_shift_rot_result[6]~q ),
	.datae(!\A_wr_data_unfiltered[0]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[6]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[6]~21 .extended_lut = "off";
defparam \A_wr_data_unfiltered[6]~21 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[6]~21 .shared_arith = "off";

dffeas \W_wr_data[6] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[6]~21_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[6]~q ),
	.prn(vcc));
defparam \W_wr_data[6] .is_wysiwyg = "true";
defparam \W_wr_data[6] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[6]~8 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[6] ),
	.datab(!\W_wr_data[6]~q ),
	.datac(!\M_alu_result[6]~q ),
	.datad(!\A_wr_data_unfiltered[6]~21_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[6]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[6]~8 .extended_lut = "off";
defparam \D_src1_reg[6]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[6]~8 .shared_arith = "off";

dffeas \E_src1[6] (
	.clk(clk_clk),
	.d(\D_src1_reg[6]~8_combout ),
	.asdata(\E_alu_result[6]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[6]~q ),
	.prn(vcc));
defparam \E_src1[6] .is_wysiwyg = "true";
defparam \E_src1[6] .power_up = "low";

cyclonev_lcell_comb \Add17~21 (
	.dataa(!\E_ctrl_alu_subtract~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!\E_src2[6]~q ),
	.datae(gnd),
	.dataf(!\E_src1[6]~q ),
	.datag(gnd),
	.cin(\Add17~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~21_sumout ),
	.cout(\Add17~22 ),
	.shareout());
defparam \Add17~21 .extended_lut = "off";
defparam \Add17~21 .lut_mask = 64'h0000FF00000055AA;
defparam \Add17~21 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result~9 (
	.dataa(!\E_src2[6]~q ),
	.datab(!\E_src1[6]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~9 .extended_lut = "off";
defparam \E_alu_result~9 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~9 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[6] (
	.dataa(!\Add17~21_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~9_combout ),
	.datae(!\E_extra_pc[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[6]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[6] .extended_lut = "off";
defparam \E_alu_result[6] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[6] .shared_arith = "off";

dffeas \M_alu_result[6] (
	.clk(clk_clk),
	.d(\E_alu_result[6]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[6]~q ),
	.prn(vcc));
defparam \M_alu_result[6] .is_wysiwyg = "true";
defparam \M_alu_result[6] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[6]~16 (
	.dataa(!\M_alu_result[6]~q ),
	.datab(!\D_src2_reg[5]~3_combout ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\W_wr_data[6]~q ),
	.datae(!\A_wr_data_unfiltered[6]~21_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[6]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[6]~16 .extended_lut = "off";
defparam \D_src2_reg[6]~16 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[6]~16 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[6]~17 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_src2_reg[6]~16_combout ),
	.datad(!\E_alu_result[6]~combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[6] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[6]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[6]~17 .extended_lut = "off";
defparam \D_src2_reg[6]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[6]~17 .shared_arith = "off";

dffeas \E_src2[6] (
	.clk(clk_clk),
	.d(\D_iw[12]~q ),
	.asdata(\D_src2_reg[6]~17_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[6]~q ),
	.prn(vcc));
defparam \E_src2[6] .is_wysiwyg = "true";
defparam \E_src2[6] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~8 (
	.dataa(!\E_src2[7]~q ),
	.datab(!\E_src1[7]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~8 .extended_lut = "off";
defparam \E_alu_result~8 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~8 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[7] (
	.dataa(!\Add17~9_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~8_combout ),
	.datae(!\E_extra_pc[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[7]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[7] .extended_lut = "off";
defparam \E_alu_result[7] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[7] .shared_arith = "off";

dffeas \M_alu_result[7] (
	.clk(clk_clk),
	.d(\E_alu_result[7]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[7]~q ),
	.prn(vcc));
defparam \M_alu_result[7] .is_wysiwyg = "true";
defparam \M_alu_result[7] .power_up = "low";

dffeas \A_inst_result[7] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.asdata(\M_alu_result[7]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[7]~q ),
	.prn(vcc));
defparam \A_inst_result[7] .is_wysiwyg = "true";
defparam \A_inst_result[7] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[7]~18 (
	.dataa(!\A_inst_result[7]~q ),
	.datab(!\A_inst_result[15]~q ),
	.datac(!\A_inst_result[23]~q ),
	.datad(!\A_inst_result[31]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[7]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[7]~18 .extended_lut = "off";
defparam \A_wr_data_unfiltered[7]~18 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[7]~18 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[7]~7 (
	.dataa(!\M_rot_prestep2[7]~q ),
	.datab(!\M_rot_prestep2[31]~q ),
	.datac(!\M_rot_prestep2[23]~q ),
	.datad(!\M_rot_prestep2[15]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~7 .extended_lut = "off";
defparam \M_rot[7]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~7 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass0~q ),
	.datac(!\M_rot_mask[7]~q ),
	.datad(!\M_rot_sel_fill0~q ),
	.datae(!\M_rot[7]~7_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~7 .extended_lut = "off";
defparam \A_shift_rot_result~7 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~7 .shared_arith = "off";

dffeas \A_shift_rot_result[7] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[7]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[7] .is_wysiwyg = "true";
defparam \A_shift_rot_result[7] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[7]~19 (
	.dataa(!\A_slow_inst_result[7]~q ),
	.datab(!\A_wr_data_unfiltered[7]~18_combout ),
	.datac(!\A_mul_result[7]~q ),
	.datad(!\A_shift_rot_result[7]~q ),
	.datae(!\A_wr_data_unfiltered[0]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[7]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[7]~19 .extended_lut = "off";
defparam \A_wr_data_unfiltered[7]~19 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[7]~19 .shared_arith = "off";

dffeas \W_wr_data[7] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[7]~19_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[7]~q ),
	.prn(vcc));
defparam \W_wr_data[7] .is_wysiwyg = "true";
defparam \W_wr_data[7] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[7]~7 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[7] ),
	.datab(!\W_wr_data[7]~q ),
	.datac(!\M_alu_result[7]~q ),
	.datad(!\A_wr_data_unfiltered[7]~19_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[7]~7 .extended_lut = "off";
defparam \D_src1_reg[7]~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[7]~7 .shared_arith = "off";

dffeas \E_src1[7] (
	.clk(clk_clk),
	.d(\D_src1_reg[7]~7_combout ),
	.asdata(\E_alu_result[7]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[7]~q ),
	.prn(vcc));
defparam \E_src1[7] .is_wysiwyg = "true";
defparam \E_src1[7] .power_up = "low";

cyclonev_lcell_comb \E_rot_step1[7]~24 (
	.dataa(!\E_src1[7]~q ),
	.datab(!\E_src1[6]~q ),
	.datac(!\E_src1[5]~q ),
	.datad(!\E_src1[4]~q ),
	.datae(!\E_src2[0]~q ),
	.dataf(!\Add7~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_step1[7]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_step1[7]~24 .extended_lut = "off";
defparam \E_rot_step1[7]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \E_rot_step1[7]~24 .shared_arith = "off";

dffeas \M_rot_prestep2[11] (
	.clk(clk_clk),
	.d(\E_rot_step1[7]~24_combout ),
	.asdata(\E_rot_step1[11]~25_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Add7~1_combout ),
	.ena(\A_stall~combout ),
	.q(\M_rot_prestep2[11]~q ),
	.prn(vcc));
defparam \M_rot_prestep2[11] .is_wysiwyg = "true";
defparam \M_rot_prestep2[11] .power_up = "low";

cyclonev_lcell_comb \M_rot[3]~3 (
	.dataa(!\M_rot_prestep2[11]~q ),
	.datab(!\M_rot_prestep2[3]~q ),
	.datac(!\M_rot_prestep2[27]~q ),
	.datad(!\M_rot_prestep2[19]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~3 .extended_lut = "off";
defparam \M_rot[3]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~3 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_sel_fill1~q ),
	.datad(!\M_rot_mask[3]~q ),
	.datae(!\M_rot[3]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~3 .extended_lut = "off";
defparam \A_shift_rot_result~3 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~3 .shared_arith = "off";

dffeas \A_shift_rot_result[11] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[11]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[11] .is_wysiwyg = "true";
defparam \A_shift_rot_result[11] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte1_data_aligned_nxt[3]~2 (
	.dataa(!\A_ld_align_sh16~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!\d_readdata_d1[27]~q ),
	.datae(!\d_readdata_d1[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte1_data_aligned_nxt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte1_data_aligned_nxt[3]~2 .extended_lut = "off";
defparam \A_slow_ld_byte1_data_aligned_nxt[3]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_slow_ld_byte1_data_aligned_nxt[3]~2 .shared_arith = "off";

dffeas \A_slow_inst_result[11] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte1_data_aligned_nxt[3]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[11]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[11] .is_wysiwyg = "true";
defparam \A_slow_inst_result[11] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[11]~10 (
	.dataa(!\A_inst_result[11]~q ),
	.datab(!\A_inst_result[27]~q ),
	.datac(!\A_slow_inst_result[11]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[11]~4_combout ),
	.dataf(!\A_wr_data_unfiltered[11]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[11]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[11]~10 .extended_lut = "off";
defparam \A_wr_data_unfiltered[11]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[11]~10 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[11]~11 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[11]~q ),
	.datad(!\A_shift_rot_result[11]~q ),
	.datae(!\A_wr_data_unfiltered[11]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[11]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[11]~11 .extended_lut = "off";
defparam \A_wr_data_unfiltered[11]~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[11]~11 .shared_arith = "off";

dffeas \W_wr_data[11] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[11]~11_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[11]~q ),
	.prn(vcc));
defparam \W_wr_data[11] .is_wysiwyg = "true";
defparam \W_wr_data[11] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[11]~10 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\A_mul_result[11]~q ),
	.datae(!\A_shift_rot_result[11]~q ),
	.dataf(!\A_wr_data_unfiltered[11]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[11]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[11]~10 .extended_lut = "off";
defparam \D_src2_reg[11]~10 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[11]~10 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[11]~94 (
	.dataa(!\M_alu_result[11]~q ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[5]~3_combout ),
	.datad(!\D_src2_reg[13]~8_combout ),
	.datae(!\W_wr_data[11]~q ),
	.dataf(!\D_src2_reg[11]~10_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[11]~94_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[11]~94 .extended_lut = "off";
defparam \D_src2_reg[11]~94 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[11]~94 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[11]~2 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[11]~q ),
	.datad(!\E_src1[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[11]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[11]~2 .extended_lut = "off";
defparam \E_logic_result[11]~2 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[11]~2 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[11]~4 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[11]~2_combout ),
	.datad(!\E_extra_pc[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[11]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[11]~4 .extended_lut = "off";
defparam \E_alu_result[11]~4 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[11]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[11]~120 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[11] ),
	.datad(!\D_src2_reg[11]~94_combout ),
	.datae(!\D_src2_reg[5]~2_combout ),
	.dataf(!\E_alu_result[11]~4_combout ),
	.datag(!\Add17~49_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[11]~120_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[11]~120 .extended_lut = "on";
defparam \D_src2_reg[11]~120 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[11]~120 .shared_arith = "off";

dffeas \E_src2[11] (
	.clk(clk_clk),
	.d(\D_iw[17]~q ),
	.asdata(\D_src2_reg[11]~120_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[11]~q ),
	.prn(vcc));
defparam \E_src2[11] .is_wysiwyg = "true";
defparam \E_src2[11] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[11] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add17~49_sumout ),
	.datac(!\E_alu_result[11]~4_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[11]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[11] .extended_lut = "off";
defparam \E_alu_result[11] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[11] .shared_arith = "off";

dffeas \M_alu_result[11] (
	.clk(clk_clk),
	.d(\E_alu_result[11]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[11]~q ),
	.prn(vcc));
defparam \M_alu_result[11] .is_wysiwyg = "true";
defparam \M_alu_result[11] .power_up = "low";

dffeas \A_inst_result[11] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[11] ),
	.asdata(\M_alu_result[11]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[11]~q ),
	.prn(vcc));
defparam \A_inst_result[11] .is_wysiwyg = "true";
defparam \A_inst_result[11] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[3]~26 (
	.dataa(!\A_inst_result[3]~q ),
	.datab(!\A_inst_result[11]~q ),
	.datac(!\A_inst_result[19]~q ),
	.datad(!\A_inst_result[27]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[3]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[3]~26 .extended_lut = "off";
defparam \A_wr_data_unfiltered[3]~26 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[3]~26 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[3]~11 (
	.dataa(!\M_rot_prestep2[3]~q ),
	.datab(!\M_rot_prestep2[27]~q ),
	.datac(!\M_rot_prestep2[19]~q ),
	.datad(!\M_rot_prestep2[11]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~11 .extended_lut = "off";
defparam \M_rot[3]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~11 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~11 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[3]~q ),
	.datac(!\M_rot_pass0~q ),
	.datad(!\M_rot_sel_fill0~q ),
	.datae(!\M_rot[3]~11_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~11 .extended_lut = "off";
defparam \A_shift_rot_result~11 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~11 .shared_arith = "off";

dffeas \A_shift_rot_result[3] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~11_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[3]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[3] .is_wysiwyg = "true";
defparam \A_shift_rot_result[3] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[3]~27 (
	.dataa(!\A_slow_inst_result[3]~q ),
	.datab(!\A_wr_data_unfiltered[3]~26_combout ),
	.datac(!\A_mul_result[3]~q ),
	.datad(!\A_shift_rot_result[3]~q ),
	.datae(!\A_wr_data_unfiltered[0]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[3]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[3]~27 .extended_lut = "off";
defparam \A_wr_data_unfiltered[3]~27 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[3]~27 .shared_arith = "off";

dffeas \W_wr_data[3] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[3]~27_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[3]~q ),
	.prn(vcc));
defparam \W_wr_data[3] .is_wysiwyg = "true";
defparam \W_wr_data[3] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[3]~11 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[3] ),
	.datab(!\W_wr_data[3]~q ),
	.datac(!\M_alu_result[3]~q ),
	.datad(!\A_wr_data_unfiltered[3]~27_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[3]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[3]~11 .extended_lut = "off";
defparam \D_src1_reg[3]~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[3]~11 .shared_arith = "off";

dffeas \E_src1[3] (
	.clk(clk_clk),
	.d(\D_src1_reg[3]~11_combout ),
	.asdata(\E_alu_result[3]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[3]~q ),
	.prn(vcc));
defparam \E_src1[3] .is_wysiwyg = "true";
defparam \E_src1[3] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~12 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src1[3]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~12 .extended_lut = "off";
defparam \E_alu_result~12 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~12 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[3] (
	.dataa(!\Add17~29_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~12_combout ),
	.datae(!\E_extra_pc[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[3]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[3] .extended_lut = "off";
defparam \E_alu_result[3] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[3] .shared_arith = "off";

dffeas \M_alu_result[3] (
	.clk(clk_clk),
	.d(\E_alu_result[3]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[3]~q ),
	.prn(vcc));
defparam \M_alu_result[3] .is_wysiwyg = "true";
defparam \M_alu_result[3] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[3]~22 (
	.dataa(!\M_alu_result[3]~q ),
	.datab(!\D_src2_reg[5]~3_combout ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\W_wr_data[3]~q ),
	.datae(!\A_wr_data_unfiltered[3]~27_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[3]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[3]~22 .extended_lut = "off";
defparam \D_src2_reg[3]~22 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[3]~22 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[3]~23 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_src2_reg[3]~22_combout ),
	.datad(!\E_alu_result[3]~combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[3] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[3]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[3]~23 .extended_lut = "off";
defparam \D_src2_reg[3]~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[3]~23 .shared_arith = "off";

dffeas \E_src2[3] (
	.clk(clk_clk),
	.d(\D_iw[9]~q ),
	.asdata(\D_src2_reg[3]~23_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[3]~q ),
	.prn(vcc));
defparam \E_src2[3] .is_wysiwyg = "true";
defparam \E_src2[3] .power_up = "low";

cyclonev_lcell_comb \E_rot_pass1~0 (
	.dataa(!\E_src2[3]~q ),
	.datab(!\E_src2[4]~q ),
	.datac(!\E_ctrl_rot~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(!\E_ctrl_shift_rot_left~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_pass1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_pass1~0 .extended_lut = "off";
defparam \E_rot_pass1~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \E_rot_pass1~0 .shared_arith = "off";

dffeas M_rot_pass1(
	.clk(clk_clk),
	.d(\E_rot_pass1~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_pass1~q ),
	.prn(vcc));
defparam M_rot_pass1.is_wysiwyg = "true";
defparam M_rot_pass1.power_up = "low";

cyclonev_lcell_comb \M_rot[4]~2 (
	.dataa(!\M_rot_prestep2[12]~q ),
	.datab(!\M_rot_prestep2[4]~q ),
	.datac(!\M_rot_prestep2[28]~q ),
	.datad(!\M_rot_prestep2[20]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~2 .extended_lut = "off";
defparam \M_rot[4]~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~2 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~2 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_pass1~q ),
	.datac(!\M_rot_sel_fill1~q ),
	.datad(!\M_rot_mask[4]~q ),
	.datae(!\M_rot[4]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~2 .extended_lut = "off";
defparam \A_shift_rot_result~2 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~2 .shared_arith = "off";

dffeas \A_shift_rot_result[12] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[12]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[12] .is_wysiwyg = "true";
defparam \A_shift_rot_result[12] .power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte1_data_aligned_nxt[4]~1 (
	.dataa(!\A_ld_align_sh16~q ),
	.datab(!\A_ld_align_byte1_fill~q ),
	.datac(!\A_slow_ld_data_fill_bit~0_combout ),
	.datad(!\d_readdata_d1[28]~q ),
	.datae(!\d_readdata_d1[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte1_data_aligned_nxt[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte1_data_aligned_nxt[4]~1 .extended_lut = "off";
defparam \A_slow_ld_byte1_data_aligned_nxt[4]~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_slow_ld_byte1_data_aligned_nxt[4]~1 .shared_arith = "off";

dffeas \A_slow_inst_result[12] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte1_data_aligned_nxt[4]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[12]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[12] .is_wysiwyg = "true";
defparam \A_slow_inst_result[12] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[12]~8 (
	.dataa(!\A_inst_result[12]~q ),
	.datab(!\A_inst_result[28]~q ),
	.datac(!\A_slow_inst_result[12]~q ),
	.datad(!\A_data_ram_ld_align_fill_bit~combout ),
	.datae(!\A_wr_data_unfiltered[11]~4_combout ),
	.dataf(!\A_wr_data_unfiltered[11]~5_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[12]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[12]~8 .extended_lut = "off";
defparam \A_wr_data_unfiltered[12]~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[12]~8 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[12]~9 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\A_mul_result[12]~q ),
	.datad(!\A_shift_rot_result[12]~q ),
	.datae(!\A_wr_data_unfiltered[12]~8_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[12]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[12]~9 .extended_lut = "off";
defparam \A_wr_data_unfiltered[12]~9 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \A_wr_data_unfiltered[12]~9 .shared_arith = "off";

dffeas \W_wr_data[12] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[12]~9_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[12]~q ),
	.prn(vcc));
defparam \W_wr_data[12] .is_wysiwyg = "true";
defparam \W_wr_data[12] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[12]~9 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_ctrl_shift_rot~q ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\A_mul_result[12]~q ),
	.datae(!\A_shift_rot_result[12]~q ),
	.dataf(!\A_wr_data_unfiltered[12]~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[12]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[12]~9 .extended_lut = "off";
defparam \D_src2_reg[12]~9 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[12]~9 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[12]~93 (
	.dataa(!\M_alu_result[12]~q ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[5]~3_combout ),
	.datad(!\D_src2_reg[13]~8_combout ),
	.datae(!\W_wr_data[12]~q ),
	.dataf(!\D_src2_reg[12]~9_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[12]~93_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[12]~93 .extended_lut = "off";
defparam \D_src2_reg[12]~93 .lut_mask = 64'hC5FFFFFFFFFFFFFF;
defparam \D_src2_reg[12]~93 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[12]~1 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[12]~q ),
	.datad(!\E_src1[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[12]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[12]~1 .extended_lut = "off";
defparam \E_logic_result[12]~1 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[12]~1 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[12]~3 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_logic_result[12]~1_combout ),
	.datad(!\E_extra_pc[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[12]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[12]~3 .extended_lut = "off";
defparam \E_alu_result[12]~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_alu_result[12]~3 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[12]~124 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[12] ),
	.datad(!\D_src2_reg[12]~93_combout ),
	.datae(!\D_src2_reg[5]~2_combout ),
	.dataf(!\E_alu_result[12]~3_combout ),
	.datag(!\Add17~45_sumout ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[12]~124_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[12]~124 .extended_lut = "on";
defparam \D_src2_reg[12]~124 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \D_src2_reg[12]~124 .shared_arith = "off";

dffeas \E_src2[12] (
	.clk(clk_clk),
	.d(\D_iw[18]~q ),
	.asdata(\D_src2_reg[12]~124_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[12]~q ),
	.prn(vcc));
defparam \E_src2[12] .is_wysiwyg = "true";
defparam \E_src2[12] .power_up = "low";

cyclonev_lcell_comb \E_alu_result[12] (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add17~45_sumout ),
	.datac(!\E_alu_result[12]~3_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[12]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[12] .extended_lut = "off";
defparam \E_alu_result[12] .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \E_alu_result[12] .shared_arith = "off";

dffeas \M_alu_result[12] (
	.clk(clk_clk),
	.d(\E_alu_result[12]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[12]~q ),
	.prn(vcc));
defparam \M_alu_result[12] .is_wysiwyg = "true";
defparam \M_alu_result[12] .power_up = "low";

dffeas \A_inst_result[12] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[12] ),
	.asdata(\M_alu_result[12]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[12]~q ),
	.prn(vcc));
defparam \A_inst_result[12] .is_wysiwyg = "true";
defparam \A_inst_result[12] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[4]~24 (
	.dataa(!\A_inst_result[4]~q ),
	.datab(!\A_inst_result[12]~q ),
	.datac(!\A_inst_result[20]~q ),
	.datad(!\A_inst_result[28]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[4]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[4]~24 .extended_lut = "off";
defparam \A_wr_data_unfiltered[4]~24 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[4]~24 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[4]~10 (
	.dataa(!\M_rot_prestep2[4]~q ),
	.datab(!\M_rot_prestep2[28]~q ),
	.datac(!\M_rot_prestep2[20]~q ),
	.datad(!\M_rot_prestep2[12]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[4]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[4]~10 .extended_lut = "off";
defparam \M_rot[4]~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[4]~10 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~10 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[4]~q ),
	.datac(!\M_rot_pass0~q ),
	.datad(!\M_rot_sel_fill0~q ),
	.datae(!\M_rot[4]~10_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~10 .extended_lut = "off";
defparam \A_shift_rot_result~10 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~10 .shared_arith = "off";

dffeas \A_shift_rot_result[4] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~10_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[4]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[4] .is_wysiwyg = "true";
defparam \A_shift_rot_result[4] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[4]~25 (
	.dataa(!\A_slow_inst_result[4]~q ),
	.datab(!\A_wr_data_unfiltered[4]~24_combout ),
	.datac(!\A_mul_result[4]~q ),
	.datad(!\A_shift_rot_result[4]~q ),
	.datae(!\A_wr_data_unfiltered[0]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[4]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[4]~25 .extended_lut = "off";
defparam \A_wr_data_unfiltered[4]~25 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[4]~25 .shared_arith = "off";

dffeas \W_wr_data[4] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[4]~25_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[4]~q ),
	.prn(vcc));
defparam \W_wr_data[4] .is_wysiwyg = "true";
defparam \W_wr_data[4] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[4]~20 (
	.dataa(!\M_alu_result[4]~q ),
	.datab(!\D_src2_reg[5]~3_combout ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\W_wr_data[4]~q ),
	.datae(!\A_wr_data_unfiltered[4]~25_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[4]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[4]~20 .extended_lut = "off";
defparam \D_src2_reg[4]~20 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[4]~20 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[4]~21 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_src2_reg[4]~20_combout ),
	.datad(!\E_alu_result[4]~combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[4] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[4]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[4]~21 .extended_lut = "off";
defparam \D_src2_reg[4]~21 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[4]~21 .shared_arith = "off";

dffeas \E_src2[4] (
	.clk(clk_clk),
	.d(\D_iw[10]~q ),
	.asdata(\D_src2_reg[4]~21_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[4]~q ),
	.prn(vcc));
defparam \E_src2[4] .is_wysiwyg = "true";
defparam \E_src2[4] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~11 (
	.dataa(!\E_src2[4]~q ),
	.datab(!\E_src1[4]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~11 .extended_lut = "off";
defparam \E_alu_result~11 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~11 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[4] (
	.dataa(!\Add17~33_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~11_combout ),
	.datae(!\E_extra_pc[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[4]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[4] .extended_lut = "off";
defparam \E_alu_result[4] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[4] .shared_arith = "off";

dffeas \M_alu_result[4] (
	.clk(clk_clk),
	.d(\E_alu_result[4]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[4]~q ),
	.prn(vcc));
defparam \M_alu_result[4] .is_wysiwyg = "true";
defparam \M_alu_result[4] .power_up = "low";

dffeas \A_mem_baddr[4] (
	.clk(clk_clk),
	.d(\M_alu_result[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[4]~q ),
	.prn(vcc));
defparam \A_mem_baddr[4] .is_wysiwyg = "true";
defparam \A_mem_baddr[4] .power_up = "low";

cyclonev_lcell_comb \A_dc_fill_has_started_nxt~0 (
	.dataa(!\A_dc_fill_has_started~q ),
	.datab(!\A_dc_fill_starting~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_has_started_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_has_started_nxt~0 .extended_lut = "off";
defparam \A_dc_fill_has_started_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \A_dc_fill_has_started_nxt~0 .shared_arith = "off";

dffeas A_dc_fill_has_started(
	.clk(clk_clk),
	.d(\A_dc_fill_has_started_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_fill_has_started~q ),
	.prn(vcc));
defparam A_dc_fill_has_started.is_wysiwyg = "true";
defparam A_dc_fill_has_started.power_up = "low";

cyclonev_lcell_comb \A_dc_fill_starting~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_want_fill~q ),
	.datac(!\A_dc_fill_has_started~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_starting~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_starting~0 .extended_lut = "off";
defparam \A_dc_fill_starting~0 .lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam \A_dc_fill_starting~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_fill_dp_offset_nxt[0]~1 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\A_dc_fill_dp_offset[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_dp_offset_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_dp_offset_nxt[0]~1 .extended_lut = "off";
defparam \A_dc_fill_dp_offset_nxt[0]~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_dc_fill_dp_offset_nxt[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_rd_data_cnt[0]~1 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_want_fill~q ),
	.datac(!\A_dc_fill_has_started~q ),
	.datad(!\d_readdatavalid_d1~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt[0]~1 .extended_lut = "off";
defparam \A_dc_rd_data_cnt[0]~1 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \A_dc_rd_data_cnt[0]~1 .shared_arith = "off";

dffeas \A_dc_fill_dp_offset[0] (
	.clk(clk_clk),
	.d(\A_dc_fill_dp_offset_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~1_combout ),
	.q(\A_dc_fill_dp_offset[0]~q ),
	.prn(vcc));
defparam \A_dc_fill_dp_offset[0] .is_wysiwyg = "true";
defparam \A_dc_fill_dp_offset[0] .power_up = "low";

cyclonev_lcell_comb \A_dc_fill_dp_offset_nxt[1]~2 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\A_dc_fill_dp_offset[0]~q ),
	.datac(!\A_dc_fill_dp_offset[1]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_dp_offset_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_dp_offset_nxt[1]~2 .extended_lut = "off";
defparam \A_dc_fill_dp_offset_nxt[1]~2 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \A_dc_fill_dp_offset_nxt[1]~2 .shared_arith = "off";

dffeas \A_dc_fill_dp_offset[1] (
	.clk(clk_clk),
	.d(\A_dc_fill_dp_offset_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~1_combout ),
	.q(\A_dc_fill_dp_offset[1]~q ),
	.prn(vcc));
defparam \A_dc_fill_dp_offset[1] .is_wysiwyg = "true";
defparam \A_dc_fill_dp_offset[1] .power_up = "low";

cyclonev_lcell_comb \A_dc_fill_dp_offset_nxt[2]~0 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\A_dc_fill_dp_offset[0]~q ),
	.datac(!\A_dc_fill_dp_offset[1]~q ),
	.datad(!\A_dc_fill_dp_offset[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_dp_offset_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_dp_offset_nxt[2]~0 .extended_lut = "off";
defparam \A_dc_fill_dp_offset_nxt[2]~0 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \A_dc_fill_dp_offset_nxt[2]~0 .shared_arith = "off";

dffeas \A_dc_fill_dp_offset[2] (
	.clk(clk_clk),
	.d(\A_dc_fill_dp_offset_nxt[2]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~1_combout ),
	.q(\A_dc_fill_dp_offset[2]~q ),
	.prn(vcc));
defparam \A_dc_fill_dp_offset[2] .is_wysiwyg = "true";
defparam \A_dc_fill_dp_offset[2] .power_up = "low";

cyclonev_lcell_comb \Equal264~0 (
	.dataa(!\A_mem_baddr[4]~q ),
	.datab(!\A_dc_fill_dp_offset[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal264~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal264~0 .extended_lut = "off";
defparam \Equal264~0 .lut_mask = 64'h6666666666666666;
defparam \Equal264~0 .shared_arith = "off";

cyclonev_lcell_comb \M_ctrl_ld_st_nxt~0 (
	.dataa(!\E_iw[1]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ctrl_ld_st_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ctrl_ld_st_nxt~0 .extended_lut = "off";
defparam \M_ctrl_ld_st_nxt~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \M_ctrl_ld_st_nxt~0 .shared_arith = "off";

dffeas M_ctrl_ld_st(
	.clk(clk_clk),
	.d(\M_ctrl_ld_st_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(!\E_iw[0]~q ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_st~q ),
	.prn(vcc));
defparam M_ctrl_ld_st.is_wysiwyg = "true";
defparam M_ctrl_ld_st.power_up = "low";

cyclonev_lcell_comb \M_valid_mem_d1~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_ld_st~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_valid_mem_d1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_valid_mem_d1~0 .extended_lut = "off";
defparam \M_valid_mem_d1~0 .lut_mask = 64'h7777777777777777;
defparam \M_valid_mem_d1~0 .shared_arith = "off";

dffeas M_valid_mem_d1(
	.clk(clk_clk),
	.d(\M_valid_mem_d1~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_valid_mem_d1~q ),
	.prn(vcc));
defparam M_valid_mem_d1.is_wysiwyg = "true";
defparam M_valid_mem_d1.power_up = "low";

dffeas \A_mem_baddr[10] (
	.clk(clk_clk),
	.d(\M_alu_result[10]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[10]~q ),
	.prn(vcc));
defparam \A_mem_baddr[10] .is_wysiwyg = "true";
defparam \A_mem_baddr[10] .power_up = "low";

dffeas \A_mem_baddr[7] (
	.clk(clk_clk),
	.d(\M_alu_result[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[7]~q ),
	.prn(vcc));
defparam \A_mem_baddr[7] .is_wysiwyg = "true";
defparam \A_mem_baddr[7] .power_up = "low";

dffeas \A_mem_baddr[6] (
	.clk(clk_clk),
	.d(\M_alu_result[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[6]~q ),
	.prn(vcc));
defparam \A_mem_baddr[6] .is_wysiwyg = "true";
defparam \A_mem_baddr[6] .power_up = "low";

dffeas \A_mem_baddr[5] (
	.clk(clk_clk),
	.d(\M_alu_result[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[5]~q ),
	.prn(vcc));
defparam \A_mem_baddr[5] .is_wysiwyg = "true";
defparam \A_mem_baddr[5] .power_up = "low";

cyclonev_lcell_comb \Equal262~0 (
	.dataa(!\A_mem_baddr[6]~q ),
	.datab(!\M_alu_result[6]~q ),
	.datac(!\A_mem_baddr[5]~q ),
	.datad(!\M_alu_result[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal262~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal262~0 .extended_lut = "off";
defparam \Equal262~0 .lut_mask = 64'h6996699669966996;
defparam \Equal262~0 .shared_arith = "off";

dffeas \A_mem_baddr[9] (
	.clk(clk_clk),
	.d(\M_alu_result[9]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[9]~q ),
	.prn(vcc));
defparam \A_mem_baddr[9] .is_wysiwyg = "true";
defparam \A_mem_baddr[9] .power_up = "low";

dffeas \A_mem_baddr[8] (
	.clk(clk_clk),
	.d(\M_alu_result[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[8]~q ),
	.prn(vcc));
defparam \A_mem_baddr[8] .is_wysiwyg = "true";
defparam \A_mem_baddr[8] .power_up = "low";

cyclonev_lcell_comb \Equal262~1 (
	.dataa(!\A_mem_baddr[9]~q ),
	.datab(!\M_alu_result[9]~q ),
	.datac(!\A_mem_baddr[8]~q ),
	.datad(!\M_alu_result[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal262~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal262~1 .extended_lut = "off";
defparam \Equal262~1 .lut_mask = 64'h6996699669966996;
defparam \Equal262~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal262~2 (
	.dataa(!\A_mem_baddr[10]~q ),
	.datab(!\M_alu_result[10]~q ),
	.datac(!\A_mem_baddr[7]~q ),
	.datad(!\M_alu_result[7]~q ),
	.datae(!\Equal262~0_combout ),
	.dataf(!\Equal262~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal262~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal262~2 .extended_lut = "off";
defparam \Equal262~2 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \Equal262~2 .shared_arith = "off";

dffeas M_A_dc_line_match_d1(
	.clk(clk_clk),
	.d(\Equal262~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\M_A_dc_line_match_d1~q ),
	.prn(vcc));
defparam M_A_dc_line_match_d1.is_wysiwyg = "true";
defparam M_A_dc_line_match_d1.power_up = "low";

cyclonev_lcell_comb A_dc_fill_need_extra_stall_nxt(
	.dataa(!\M_alu_result[4]~q ),
	.datab(!\M_alu_result[3]~q ),
	.datac(!\M_alu_result[2]~q ),
	.datad(!\M_valid_mem_d1~q ),
	.datae(!\M_A_dc_line_match_d1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_need_extra_stall_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_fill_need_extra_stall_nxt.extended_lut = "off";
defparam A_dc_fill_need_extra_stall_nxt.lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam A_dc_fill_need_extra_stall_nxt.shared_arith = "off";

dffeas A_dc_fill_need_extra_stall(
	.clk(clk_clk),
	.d(\A_dc_fill_need_extra_stall_nxt~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_fill_need_extra_stall~q ),
	.prn(vcc));
defparam A_dc_fill_need_extra_stall.is_wysiwyg = "true";
defparam A_dc_fill_need_extra_stall.power_up = "low";

cyclonev_lcell_comb \A_dc_rd_data_cnt_nxt[0]~3 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\d_readdatavalid_d1~q ),
	.datac(!\A_dc_rd_data_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt_nxt[0]~3 .extended_lut = "off";
defparam \A_dc_rd_data_cnt_nxt[0]~3 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \A_dc_rd_data_cnt_nxt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_rd_data_cnt[0]~0 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_dc_wb_active~q ),
	.datac(!\A_dc_want_fill~q ),
	.datad(!\A_dc_fill_has_started~q ),
	.datae(!\d_readdatavalid_d1~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt[0]~0 .extended_lut = "off";
defparam \A_dc_rd_data_cnt[0]~0 .lut_mask = 64'hFFEFFFFFFFEFFFFF;
defparam \A_dc_rd_data_cnt[0]~0 .shared_arith = "off";

dffeas \A_dc_rd_data_cnt[0] (
	.clk(clk_clk),
	.d(\A_dc_rd_data_cnt_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~0_combout ),
	.q(\A_dc_rd_data_cnt[0]~q ),
	.prn(vcc));
defparam \A_dc_rd_data_cnt[0] .is_wysiwyg = "true";
defparam \A_dc_rd_data_cnt[0] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_data_cnt_nxt[1]~2 (
	.dataa(!\d_readdatavalid_d1~q ),
	.datab(!\A_dc_rd_data_cnt[1]~q ),
	.datac(!\A_dc_rd_data_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt_nxt[1]~2 .extended_lut = "off";
defparam \A_dc_rd_data_cnt_nxt[1]~2 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \A_dc_rd_data_cnt_nxt[1]~2 .shared_arith = "off";

dffeas \A_dc_rd_data_cnt[1] (
	.clk(clk_clk),
	.d(\A_dc_rd_data_cnt_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~0_combout ),
	.q(\A_dc_rd_data_cnt[1]~q ),
	.prn(vcc));
defparam \A_dc_rd_data_cnt[1] .is_wysiwyg = "true";
defparam \A_dc_rd_data_cnt[1] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_data_cnt_nxt[2]~1 (
	.dataa(!\d_readdatavalid_d1~q ),
	.datab(!\A_dc_rd_data_cnt[2]~q ),
	.datac(!\A_dc_rd_data_cnt[1]~q ),
	.datad(!\A_dc_rd_data_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt_nxt[2]~1 .extended_lut = "off";
defparam \A_dc_rd_data_cnt_nxt[2]~1 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \A_dc_rd_data_cnt_nxt[2]~1 .shared_arith = "off";

dffeas \A_dc_rd_data_cnt[2] (
	.clk(clk_clk),
	.d(\A_dc_rd_data_cnt_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~0_combout ),
	.q(\A_dc_rd_data_cnt[2]~q ),
	.prn(vcc));
defparam \A_dc_rd_data_cnt[2] .is_wysiwyg = "true";
defparam \A_dc_rd_data_cnt[2] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_data_cnt_nxt[3]~0 (
	.dataa(!\A_dc_fill_starting~0_combout ),
	.datab(!\A_dc_rd_data_cnt[3]~q ),
	.datac(!\d_readdatavalid_d1~q ),
	.datad(!\A_dc_rd_data_cnt[2]~q ),
	.datae(!\A_dc_rd_data_cnt[1]~q ),
	.dataf(!\A_dc_rd_data_cnt[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_data_cnt_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_data_cnt_nxt[3]~0 .extended_lut = "off";
defparam \A_dc_rd_data_cnt_nxt[3]~0 .lut_mask = 64'hEBBEBEEBBEEBEBBE;
defparam \A_dc_rd_data_cnt_nxt[3]~0 .shared_arith = "off";

dffeas \A_dc_rd_data_cnt[3] (
	.clk(clk_clk),
	.d(\A_dc_rd_data_cnt_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_data_cnt[0]~0_combout ),
	.q(\A_dc_rd_data_cnt[3]~q ),
	.prn(vcc));
defparam \A_dc_rd_data_cnt[3] .is_wysiwyg = "true";
defparam \A_dc_rd_data_cnt[3] .power_up = "low";

cyclonev_lcell_comb A_ld_bypass_done(
	.dataa(!\A_dc_rd_data_cnt[3]~q ),
	.datab(!\d_readdatavalid_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_ld_bypass_done~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_ld_bypass_done.extended_lut = "off";
defparam A_ld_bypass_done.lut_mask = 64'h7777777777777777;
defparam A_ld_bypass_done.shared_arith = "off";

dffeas A_dc_rd_last_transfer_d1(
	.clk(clk_clk),
	.d(\A_ld_bypass_done~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_rd_last_transfer_d1~q ),
	.prn(vcc));
defparam A_dc_rd_last_transfer_d1.is_wysiwyg = "true";
defparam A_dc_rd_last_transfer_d1.power_up = "low";

cyclonev_lcell_comb \A_dc_fill_active_nxt~0 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_dc_fill_starting~0_combout ),
	.datac(!\A_dc_fill_need_extra_stall~q ),
	.datad(!\A_dc_rd_last_transfer_d1~q ),
	.datae(!\A_ld_bypass_done~combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_active_nxt~0 .extended_lut = "off";
defparam \A_dc_fill_active_nxt~0 .lut_mask = 64'hFFFFFF7BFFFFFF7B;
defparam \A_dc_fill_active_nxt~0 .shared_arith = "off";

dffeas A_dc_fill_active(
	.clk(clk_clk),
	.d(\A_dc_fill_active_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_fill_active~q ),
	.prn(vcc));
defparam A_dc_fill_active.is_wysiwyg = "true";
defparam A_dc_fill_active.power_up = "low";

dffeas \A_mem_baddr[3] (
	.clk(clk_clk),
	.d(\M_alu_result[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[3]~q ),
	.prn(vcc));
defparam \A_mem_baddr[3] .is_wysiwyg = "true";
defparam \A_mem_baddr[3] .power_up = "low";

dffeas \A_mem_baddr[2] (
	.clk(clk_clk),
	.d(\M_alu_result[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[2]~q ),
	.prn(vcc));
defparam \A_mem_baddr[2] .is_wysiwyg = "true";
defparam \A_mem_baddr[2] .power_up = "low";

cyclonev_lcell_comb \A_dc_fill_wr_data~0 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_mem_baddr[3]~q ),
	.datac(!\A_mem_baddr[2]~q ),
	.datad(!\A_dc_fill_dp_offset[0]~q ),
	.datae(!\A_dc_fill_dp_offset[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_fill_wr_data~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_fill_wr_data~0 .extended_lut = "off";
defparam \A_dc_fill_wr_data~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \A_dc_fill_wr_data~0 .shared_arith = "off";

cyclonev_lcell_comb \A_slow_inst_result_en~0 (
	.dataa(!\d_readdatavalid_d1~q ),
	.datab(!\A_ctrl_ld_bypass~q ),
	.datac(!\Equal264~0_combout ),
	.datad(!\A_dc_fill_wr_data~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_inst_result_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_inst_result_en~0 .extended_lut = "off";
defparam \A_slow_inst_result_en~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \A_slow_inst_result_en~0 .shared_arith = "off";

dffeas \A_slow_inst_result[1] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte0_data_aligned_nxt[1]~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[1]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[1] .is_wysiwyg = "true";
defparam \A_slow_inst_result[1] .power_up = "low";

dffeas \A_inst_result[1] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(\M_alu_result[1]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[1]~q ),
	.prn(vcc));
defparam \A_inst_result[1] .is_wysiwyg = "true";
defparam \A_inst_result[1] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[1]~28 (
	.dataa(!\A_inst_result[1]~q ),
	.datab(!\A_inst_result[9]~q ),
	.datac(!\A_inst_result[17]~q ),
	.datad(!\A_inst_result[25]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[1]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[1]~28 .extended_lut = "off";
defparam \A_wr_data_unfiltered[1]~28 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[1]~28 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[1]~12 (
	.dataa(!\M_rot_prestep2[1]~q ),
	.datab(!\M_rot_prestep2[25]~q ),
	.datac(!\M_rot_prestep2[17]~q ),
	.datad(!\M_rot_prestep2[9]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[1]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[1]~12 .extended_lut = "off";
defparam \M_rot[1]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[1]~12 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~12 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[1]~q ),
	.datac(!\M_rot_pass0~q ),
	.datad(!\M_rot_sel_fill0~q ),
	.datae(!\M_rot[1]~12_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~12 .extended_lut = "off";
defparam \A_shift_rot_result~12 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~12 .shared_arith = "off";

dffeas \A_shift_rot_result[1] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~12_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[1]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[1] .is_wysiwyg = "true";
defparam \A_shift_rot_result[1] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[1]~29 (
	.dataa(!\A_slow_inst_result[1]~q ),
	.datab(!\A_wr_data_unfiltered[1]~28_combout ),
	.datac(!\A_mul_result[1]~q ),
	.datad(!\A_shift_rot_result[1]~q ),
	.datae(!\A_wr_data_unfiltered[0]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[1]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[1]~29 .extended_lut = "off";
defparam \A_wr_data_unfiltered[1]~29 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[1]~29 .shared_arith = "off";

dffeas \W_wr_data[1] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[1]~29_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[1]~q ),
	.prn(vcc));
defparam \W_wr_data[1] .is_wysiwyg = "true";
defparam \W_wr_data[1] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[1]~24 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\W_wr_data[1]~q ),
	.datad(!\A_wr_data_unfiltered[1]~29_combout ),
	.datae(!\M_alu_result[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[1]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[1]~24 .extended_lut = "off";
defparam \D_src2_reg[1]~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[1]~24 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[1]~25 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_src2_reg[1]~24_combout ),
	.datad(!\E_alu_result[1]~combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[1] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[1]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[1]~25 .extended_lut = "off";
defparam \D_src2_reg[1]~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[1]~25 .shared_arith = "off";

dffeas \E_src2[1] (
	.clk(clk_clk),
	.d(\D_iw[7]~q ),
	.asdata(\D_src2_reg[1]~25_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[1]~q ),
	.prn(vcc));
defparam \E_src2[1] .is_wysiwyg = "true";
defparam \E_src2[1] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[1]~12 (
	.dataa(!\E_src2[1]~q ),
	.datab(!\E_src1[1]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[1]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[1]~12 .extended_lut = "off";
defparam \E_logic_result[1]~12 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[1]~12 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[1] (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add17~53_sumout ),
	.datad(!\E_logic_result[1]~12_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[1]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[1] .extended_lut = "off";
defparam \E_alu_result[1] .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \E_alu_result[1] .shared_arith = "off";

dffeas \M_alu_result[1] (
	.clk(clk_clk),
	.d(\E_alu_result[1]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[1]~q ),
	.prn(vcc));
defparam \M_alu_result[1] .is_wysiwyg = "true";
defparam \M_alu_result[1] .power_up = "low";

cyclonev_lcell_comb \M_ld_align_sh16~0 (
	.dataa(!\M_alu_result[1]~q ),
	.datab(!\M_ctrl_ld8~q ),
	.datac(!\M_ctrl_ld16~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ld_align_sh16~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ld_align_sh16~0 .extended_lut = "off";
defparam \M_ld_align_sh16~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_ld_align_sh16~0 .shared_arith = "off";

dffeas A_ld_align_sh16(
	.clk(clk_clk),
	.d(\M_ld_align_sh16~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ld_align_sh16~q ),
	.prn(vcc));
defparam A_ld_align_sh16.is_wysiwyg = "true";
defparam A_ld_align_sh16.power_up = "low";

cyclonev_lcell_comb \A_slow_ld_byte0_data_aligned_nxt[2]~0 (
	.dataa(!\d_readdata_d1[2]~q ),
	.datab(!\d_readdata_d1[10]~q ),
	.datac(!\d_readdata_d1[18]~q ),
	.datad(!\d_readdata_d1[26]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_slow_ld_byte0_data_aligned_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_slow_ld_byte0_data_aligned_nxt[2]~0 .extended_lut = "off";
defparam \A_slow_ld_byte0_data_aligned_nxt[2]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_slow_ld_byte0_data_aligned_nxt[2]~0 .shared_arith = "off";

dffeas \A_slow_inst_result[2] (
	.clk(clk_clk),
	.d(\A_slow_ld_byte0_data_aligned_nxt[2]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[2]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[2] .is_wysiwyg = "true";
defparam \A_slow_inst_result[2] .power_up = "low";

dffeas \A_inst_result[2] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(\M_alu_result[2]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\M_ctrl_rdctl_inst~q ),
	.sload(!\M_ctrl_mem~q ),
	.ena(\A_stall~combout ),
	.q(\A_inst_result[2]~q ),
	.prn(vcc));
defparam \A_inst_result[2] .is_wysiwyg = "true";
defparam \A_inst_result[2] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[2]~0 (
	.dataa(!\A_inst_result[2]~q ),
	.datab(!\A_inst_result[10]~q ),
	.datac(!\A_inst_result[18]~q ),
	.datad(!\A_inst_result[26]~q ),
	.datae(!\A_ld_align_sh8~q ),
	.dataf(!\A_ld_align_sh16~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[2]~0 .extended_lut = "off";
defparam \A_wr_data_unfiltered[2]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \M_rot[2]~0 (
	.dataa(!\M_rot_prestep2[2]~q ),
	.datab(!\M_rot_prestep2[26]~q ),
	.datac(!\M_rot_prestep2[18]~q ),
	.datad(!\M_rot_prestep2[10]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[2]~0 .extended_lut = "off";
defparam \M_rot[2]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~0 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[2]~q ),
	.datac(!\M_rot_pass0~q ),
	.datad(!\M_rot_sel_fill0~q ),
	.datae(!\M_rot[2]~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~0 .extended_lut = "off";
defparam \A_shift_rot_result~0 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~0 .shared_arith = "off";

dffeas \A_shift_rot_result[2] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[2]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[2] .is_wysiwyg = "true";
defparam \A_shift_rot_result[2] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[2]~3 (
	.dataa(!\A_slow_inst_result[2]~q ),
	.datab(!\A_wr_data_unfiltered[2]~0_combout ),
	.datac(!\A_mul_result[2]~q ),
	.datad(!\A_shift_rot_result[2]~q ),
	.datae(!\A_wr_data_unfiltered[0]~1_combout ),
	.dataf(!\A_wr_data_unfiltered[0]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[2]~3 .extended_lut = "off";
defparam \A_wr_data_unfiltered[2]~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \A_wr_data_unfiltered[2]~3 .shared_arith = "off";

dffeas \W_wr_data[2] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[2]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[2]~q ),
	.prn(vcc));
defparam \W_wr_data[2] .is_wysiwyg = "true";
defparam \W_wr_data[2] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[2]~0 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[2] ),
	.datab(!\W_wr_data[2]~q ),
	.datac(!\M_alu_result[2]~q ),
	.datad(!\A_wr_data_unfiltered[2]~3_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[2]~0 .extended_lut = "off";
defparam \D_src1_reg[2]~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[2]~0 .shared_arith = "off";

dffeas \E_src1[2] (
	.clk(clk_clk),
	.d(\D_src1_reg[2]~0_combout ),
	.asdata(\E_alu_result[2]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[2]~q ),
	.prn(vcc));
defparam \E_src1[2] .is_wysiwyg = "true";
defparam \E_src1[2] .power_up = "low";

cyclonev_lcell_comb \E_alu_result~1 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src1[2]~q ),
	.datac(!\E_ctrl_logic~q ),
	.datad(!\E_logic_op[1]~q ),
	.datae(!\E_logic_op[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result~1 .extended_lut = "off";
defparam \E_alu_result~1 .lut_mask = 64'h6F9F9F6F6F9F9F6F;
defparam \E_alu_result~1 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[2] (
	.dataa(!\Add17~25_sumout ),
	.datab(!\E_ctrl_retaddr~q ),
	.datac(!\E_alu_result~0_combout ),
	.datad(!\E_alu_result~1_combout ),
	.datae(!\E_extra_pc[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[2]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[2] .extended_lut = "off";
defparam \E_alu_result[2] .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_alu_result[2] .shared_arith = "off";

dffeas \M_alu_result[2] (
	.clk(clk_clk),
	.d(\E_alu_result[2]~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_alu_result[2]~q ),
	.prn(vcc));
defparam \M_alu_result[2] .is_wysiwyg = "true";
defparam \M_alu_result[2] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[2]~5 (
	.dataa(!\M_alu_result[2]~q ),
	.datab(!\D_src2_reg[5]~3_combout ),
	.datac(!\D_src2_reg[5]~4_combout ),
	.datad(!\W_wr_data[2]~q ),
	.datae(!\A_wr_data_unfiltered[2]~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[2]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[2]~5 .extended_lut = "off";
defparam \D_src2_reg[2]~5 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \D_src2_reg[2]~5 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[2]~6 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_src2_reg[2]~5_combout ),
	.datad(!\E_alu_result[2]~combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[2] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[2]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[2]~6 .extended_lut = "off";
defparam \D_src2_reg[2]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[2]~6 .shared_arith = "off";

dffeas \E_src2[2] (
	.clk(clk_clk),
	.d(\D_iw[8]~q ),
	.asdata(\D_src2_reg[2]~6_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[2]~q ),
	.prn(vcc));
defparam \E_src2[2] .is_wysiwyg = "true";
defparam \E_src2[2] .power_up = "low";

cyclonev_lcell_comb \E_rot_mask[3]~3 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src2[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_ctrl_shift_rot_right~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_rot_mask[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_rot_mask[3]~3 .extended_lut = "off";
defparam \E_rot_mask[3]~3 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_rot_mask[3]~3 .shared_arith = "off";

dffeas \M_rot_mask[3] (
	.clk(clk_clk),
	.d(\E_rot_mask[3]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_rot_mask[3]~q ),
	.prn(vcc));
defparam \M_rot_mask[3] .is_wysiwyg = "true";
defparam \M_rot_mask[3] .power_up = "low";

cyclonev_lcell_comb \M_rot[3]~20 (
	.dataa(!\M_rot_prestep2[27]~q ),
	.datab(!\M_rot_prestep2[19]~q ),
	.datac(!\M_rot_prestep2[11]~q ),
	.datad(!\M_rot_prestep2[3]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[3]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[3]~20 .extended_lut = "off";
defparam \M_rot[3]~20 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[3]~20 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~20 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[3]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[3]~20_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~20 .extended_lut = "off";
defparam \A_shift_rot_result~20 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~20 .shared_arith = "off";

dffeas \A_shift_rot_result[27] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~20_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[27]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[27] .is_wysiwyg = "true";
defparam \A_shift_rot_result[27] .power_up = "low";

dffeas \A_slow_inst_result[27] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[27]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[27]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[27] .is_wysiwyg = "true";
defparam \A_slow_inst_result[27] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[27]~45 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[27]~q ),
	.dataf(!\A_slow_inst_result[27]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[27]~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[27]~45 .extended_lut = "off";
defparam \A_wr_data_unfiltered[27]~45 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[27]~45 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[27]~46 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[27]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[27]~q ),
	.datae(!\A_wr_data_unfiltered[27]~45_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[27]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[27]~46 .extended_lut = "off";
defparam \A_wr_data_unfiltered[27]~46 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[27]~46 .shared_arith = "off";

dffeas \W_wr_data[27] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[27]~46_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[27]~q ),
	.prn(vcc));
defparam \W_wr_data[27] .is_wysiwyg = "true";
defparam \W_wr_data[27] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[27]~12 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[27] ),
	.datab(!\W_wr_data[27]~q ),
	.datac(!\M_alu_result[27]~q ),
	.datad(!\A_wr_data_unfiltered[27]~46_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[27]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[27]~12 .extended_lut = "off";
defparam \D_src1_reg[27]~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[27]~12 .shared_arith = "off";

dffeas \E_src1[27] (
	.clk(clk_clk),
	.d(\D_src1_reg[27]~12_combout ),
	.asdata(\E_alu_result[27]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[27]~q ),
	.prn(vcc));
defparam \E_src1[27] .is_wysiwyg = "true";
defparam \E_src1[27] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[27]~56 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~20_combout ),
	.datad(!\Add17~97_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~56 .extended_lut = "off";
defparam \D_src2_reg[27]~56 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[27]~56 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~41 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[27]~q ),
	.datae(!\A_wr_data_unfiltered[27]~46_combout ),
	.dataf(!\M_alu_result[27]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~41 .extended_lut = "off";
defparam \D_src2_reg[27]~41 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[27]~41 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[27]~0 (
	.dataa(!\D_ctrl_hi_imm16~q ),
	.datab(!\D_iw[17]~q ),
	.datac(!\D_iw[21]~q ),
	.datad(!\D_ctrl_unsigned_lo_imm16~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[27]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[27]~0 .extended_lut = "off";
defparam \D_src2[27]~0 .lut_mask = 64'h7FBF7FBF7FBF7FBF;
defparam \D_src2[27]~0 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[27]~1 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[27]~56_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.datae(!\D_src2_reg[27]~41_combout ),
	.dataf(!\D_src2[27]~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[27]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[27]~1 .extended_lut = "off";
defparam \D_src2[27]~1 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[27]~1 .shared_arith = "off";

dffeas \E_src2[27] (
	.clk(clk_clk),
	.d(\D_src2[27]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[19]~1_combout ),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[27]~q ),
	.prn(vcc));
defparam \E_src2[27] .is_wysiwyg = "true";
defparam \E_src2[27] .power_up = "low";

cyclonev_lcell_comb \E_logic_result[27]~6 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[27]~q ),
	.datad(!\E_src1[27]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[27]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[27]~6 .extended_lut = "off";
defparam \E_logic_result[27]~6 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[27]~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~0 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[17]~q ),
	.datad(!\E_src1[17]~q ),
	.datae(!\E_src2[16]~q ),
	.dataf(!\E_src1[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~0 .extended_lut = "off";
defparam \Equal303~0 .lut_mask = 64'h6996966996696996;
defparam \Equal303~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~1 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[28]~q ),
	.datad(!\E_src1[28]~q ),
	.datae(!\E_src2[18]~q ),
	.dataf(!\E_src1[18]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~1 .extended_lut = "off";
defparam \Equal303~1 .lut_mask = 64'h6996966996696996;
defparam \Equal303~1 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~2 (
	.dataa(!\E_logic_result[27]~6_combout ),
	.datab(!\E_logic_result[29]~7_combout ),
	.datac(!\E_logic_result[30]~8_combout ),
	.datad(!\E_logic_result[31]~9_combout ),
	.datae(!\Equal303~0_combout ),
	.dataf(!\Equal303~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~2 .extended_lut = "off";
defparam \Equal303~2 .lut_mask = 64'hFFFEFFFFFFFFFFFF;
defparam \Equal303~2 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~3 (
	.dataa(!\E_src2[2]~q ),
	.datab(!\E_src1[2]~q ),
	.datac(!\E_src2[3]~q ),
	.datad(!\E_src1[3]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~3 .extended_lut = "off";
defparam \Equal303~3 .lut_mask = 64'h6996966996696996;
defparam \Equal303~3 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~4 (
	.dataa(!\E_src2[4]~q ),
	.datab(!\E_src1[4]~q ),
	.datac(!\E_src2[5]~q ),
	.datad(!\E_src1[5]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~4 .extended_lut = "off";
defparam \Equal303~4 .lut_mask = 64'h6996966996696996;
defparam \Equal303~4 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~5 (
	.dataa(!\E_src2[6]~q ),
	.datab(!\E_src1[6]~q ),
	.datac(!\E_src2[7]~q ),
	.datad(!\E_src1[7]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~5 .extended_lut = "off";
defparam \Equal303~5 .lut_mask = 64'h6996966996696996;
defparam \Equal303~5 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~6 (
	.dataa(!\E_src2[8]~q ),
	.datab(!\E_src1[8]~q ),
	.datac(!\E_src2[9]~q ),
	.datad(!\E_src1[9]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~6 .extended_lut = "off";
defparam \Equal303~6 .lut_mask = 64'h6996966996696996;
defparam \Equal303~6 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~7 (
	.dataa(!\E_src2[13]~q ),
	.datab(!\E_src1[13]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_src2[12]~q ),
	.dataf(!\E_src1[12]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~7 .extended_lut = "off";
defparam \Equal303~7 .lut_mask = 64'h6996966996696996;
defparam \Equal303~7 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~8 (
	.dataa(!\E_src2[10]~q ),
	.datab(!\E_src1[10]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(!\E_src2[11]~q ),
	.dataf(!\E_src1[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~8 .extended_lut = "off";
defparam \Equal303~8 .lut_mask = 64'h6996966996696996;
defparam \Equal303~8 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~9 (
	.dataa(!\Equal303~3_combout ),
	.datab(!\Equal303~4_combout ),
	.datac(!\Equal303~5_combout ),
	.datad(!\Equal303~6_combout ),
	.datae(!\Equal303~7_combout ),
	.dataf(!\Equal303~8_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~9 .extended_lut = "off";
defparam \Equal303~9 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \Equal303~9 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~10 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[26]~q ),
	.datad(!\E_src1[26]~q ),
	.datae(!\E_src2[19]~q ),
	.dataf(!\E_src1[19]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~10 .extended_lut = "off";
defparam \Equal303~10 .lut_mask = 64'h6996966996696996;
defparam \Equal303~10 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~11 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[25]~q ),
	.datad(!\E_src1[25]~q ),
	.datae(!\E_src2[20]~q ),
	.dataf(!\E_src1[20]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~11 .extended_lut = "off";
defparam \Equal303~11 .lut_mask = 64'h6996966996696996;
defparam \Equal303~11 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~12 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[22]~q ),
	.datad(!\E_src1[22]~q ),
	.datae(!\E_src2[14]~q ),
	.dataf(!\E_src1[14]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~12 .extended_lut = "off";
defparam \Equal303~12 .lut_mask = 64'h6996966996696996;
defparam \Equal303~12 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~13 (
	.dataa(!\E_logic_op[1]~q ),
	.datab(!\E_logic_op[0]~q ),
	.datac(!\E_src2[24]~q ),
	.datad(!\E_src1[24]~q ),
	.datae(!\E_src2[23]~q ),
	.dataf(!\E_src1[23]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~13 .extended_lut = "off";
defparam \Equal303~13 .lut_mask = 64'h6996966996696996;
defparam \Equal303~13 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~14 (
	.dataa(!\E_src2[1]~q ),
	.datab(!\E_src1[1]~q ),
	.datac(!\E_src2[0]~q ),
	.datad(!\E_src1[0]~q ),
	.datae(!\E_logic_op[1]~q ),
	.dataf(!\E_logic_op[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~14 .extended_lut = "off";
defparam \Equal303~14 .lut_mask = 64'h6996966996696996;
defparam \Equal303~14 .shared_arith = "off";

cyclonev_lcell_comb \Equal303~15 (
	.dataa(!\E_logic_result[21]~10_combout ),
	.datab(!\E_logic_result[15]~11_combout ),
	.datac(!\Equal303~11_combout ),
	.datad(!\Equal303~12_combout ),
	.datae(!\Equal303~13_combout ),
	.dataf(!\Equal303~14_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal303~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal303~15 .extended_lut = "off";
defparam \Equal303~15 .lut_mask = 64'hEFFFFFFFFFFFFFFF;
defparam \Equal303~15 .shared_arith = "off";

dffeas \E_compare_op[1] (
	.clk(clk_clk),
	.d(\D_logic_op_raw[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_compare_op[1]~q ),
	.prn(vcc));
defparam \E_compare_op[1] .is_wysiwyg = "true";
defparam \E_compare_op[1] .power_up = "low";

cyclonev_lcell_comb \E_br_result~0 (
	.dataa(!\E_compare_op[0]~q ),
	.datab(!\Equal303~2_combout ),
	.datac(!\Equal303~9_combout ),
	.datad(!\Equal303~10_combout ),
	.datae(!\Equal303~15_combout ),
	.dataf(!\E_compare_op[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_result~0 .extended_lut = "off";
defparam \E_br_result~0 .lut_mask = 64'hFFFFFFFF7DD7D77D;
defparam \E_br_result~0 .shared_arith = "off";

cyclonev_lcell_comb \E_br_result~1 (
	.dataa(!\E_compare_op[0]~q ),
	.datab(!\Equal303~2_combout ),
	.datac(!\Equal303~9_combout ),
	.datad(!\Equal303~10_combout ),
	.datae(!\Equal303~15_combout ),
	.dataf(!\E_compare_op[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_result~1 .extended_lut = "off";
defparam \E_br_result~1 .lut_mask = 64'hBEEBEBBEFFFFFFFF;
defparam \E_br_result~1 .shared_arith = "off";

cyclonev_lcell_comb \E_logic_result[0]~13 (
	.dataa(!\E_src2[0]~q ),
	.datab(!\E_src1[0]~q ),
	.datac(!\E_logic_op[1]~q ),
	.datad(!\E_logic_op[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_logic_result[0]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_logic_result[0]~13 .extended_lut = "off";
defparam \E_logic_result[0]~13 .lut_mask = 64'h6996699669966996;
defparam \E_logic_result[0]~13 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[0]~13 (
	.dataa(!\E_ctrl_logic~q ),
	.datab(!\E_alu_result~0_combout ),
	.datac(!\Add17~57_sumout ),
	.datad(!\E_logic_result[0]~13_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[0]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[0]~13 .extended_lut = "off";
defparam \E_alu_result[0]~13 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \E_alu_result[0]~13 .shared_arith = "off";

cyclonev_lcell_comb \E_alu_result[0] (
	.dataa(!\E_ctrl_cmp~q ),
	.datab(!\Add17~61_sumout ),
	.datac(!\E_br_result~0_combout ),
	.datad(!\E_br_result~1_combout ),
	.datae(!\E_alu_result[0]~13_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_alu_result[0]~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_alu_result[0] .extended_lut = "off";
defparam \E_alu_result[0] .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \E_alu_result[0] .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~26 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\W_wr_data[0]~q ),
	.datad(!\A_wr_data_unfiltered[0]~31_combout ),
	.datae(!\M_alu_result[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~26 .extended_lut = "off";
defparam \D_src2_reg[0]~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[0]~26 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[0]~27 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\E_alu_result[0]~combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[0] ),
	.datae(!\D_src2_reg[0]~26_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[0]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[0]~27 .extended_lut = "off";
defparam \D_src2_reg[0]~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[0]~27 .shared_arith = "off";

dffeas \E_src2[0] (
	.clk(clk_clk),
	.d(\D_iw[6]~q ),
	.asdata(\D_src2_reg[0]~27_combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\E_src2[14]~0_combout ),
	.sload(!\D_ctrl_src2_choose_imm~q ),
	.ena(\A_stall~combout ),
	.q(\E_src2[0]~q ),
	.prn(vcc));
defparam \E_src2[0] .is_wysiwyg = "true";
defparam \E_src2[0] .power_up = "low";

cyclonev_lcell_comb \M_data_ram_ld_align_sign_bit_16_hi~0 (
	.dataa(!\Add17~57_sumout ),
	.datab(!\Equal187~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_data_ram_ld_align_sign_bit_16_hi~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_data_ram_ld_align_sign_bit_16_hi~0 .extended_lut = "off";
defparam \M_data_ram_ld_align_sign_bit_16_hi~0 .lut_mask = 64'h7777777777777777;
defparam \M_data_ram_ld_align_sign_bit_16_hi~0 .shared_arith = "off";

dffeas M_data_ram_ld_align_sign_bit_16_hi(
	.clk(clk_clk),
	.d(\M_data_ram_ld_align_sign_bit_16_hi~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_data_ram_ld_align_sign_bit_16_hi~q ),
	.prn(vcc));
defparam M_data_ram_ld_align_sign_bit_16_hi.is_wysiwyg = "true";
defparam M_data_ram_ld_align_sign_bit_16_hi.power_up = "low";

cyclonev_lcell_comb \M_data_ram_ld_align_sign_bit~0 (
	.dataa(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[7] ),
	.datab(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[15] ),
	.datac(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[23] ),
	.datad(!\embedded_system_nios2_qsys_0_dc_data|the_altsyncram|auto_generated|q_b[31] ),
	.datae(!\M_data_ram_ld_align_sign_bit_16_hi~q ),
	.dataf(!\M_alu_result[1]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_data_ram_ld_align_sign_bit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_data_ram_ld_align_sign_bit~0 .extended_lut = "off";
defparam \M_data_ram_ld_align_sign_bit~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_data_ram_ld_align_sign_bit~0 .shared_arith = "off";

dffeas A_data_ram_ld_align_sign_bit(
	.clk(clk_clk),
	.d(\M_data_ram_ld_align_sign_bit~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_data_ram_ld_align_sign_bit~q ),
	.prn(vcc));
defparam A_data_ram_ld_align_sign_bit.is_wysiwyg = "true";
defparam A_data_ram_ld_align_sign_bit.power_up = "low";

cyclonev_lcell_comb \M_rot[7]~30 (
	.dataa(!\M_rot_prestep2[31]~q ),
	.datab(!\M_rot_prestep2[23]~q ),
	.datac(!\M_rot_prestep2[15]~q ),
	.datad(!\M_rot_prestep2[7]~q ),
	.datae(!\M_rot_rn[3]~q ),
	.dataf(!\M_rot_rn[4]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_rot[7]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_rot[7]~30 .extended_lut = "off";
defparam \M_rot[7]~30 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \M_rot[7]~30 .shared_arith = "off";

cyclonev_lcell_comb \A_shift_rot_result~30 (
	.dataa(!\M_rot_fill_bit~q ),
	.datab(!\M_rot_mask[7]~q ),
	.datac(!\M_rot_pass3~q ),
	.datad(!\M_rot_sel_fill3~q ),
	.datae(!\M_rot[7]~30_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_shift_rot_result~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_shift_rot_result~30 .extended_lut = "off";
defparam \A_shift_rot_result~30 .lut_mask = 64'hD77DFFFFD77DFFFF;
defparam \A_shift_rot_result~30 .shared_arith = "off";

dffeas \A_shift_rot_result[31] (
	.clk(clk_clk),
	.d(\A_shift_rot_result~30_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_shift_rot_result[31]~q ),
	.prn(vcc));
defparam \A_shift_rot_result[31] .is_wysiwyg = "true";
defparam \A_shift_rot_result[31] .power_up = "low";

dffeas \A_slow_inst_result[31] (
	.clk(clk_clk),
	.d(\A_slow_ld_data_fill_bit~0_combout ),
	.asdata(\d_readdata_d1[31]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\A_ld_align_byte2_byte3_fill~q ),
	.ena(\A_slow_inst_result_en~0_combout ),
	.q(\A_slow_inst_result[31]~q ),
	.prn(vcc));
defparam \A_slow_inst_result[31] .is_wysiwyg = "true";
defparam \A_slow_inst_result[31] .power_up = "low";

cyclonev_lcell_comb \A_wr_data_unfiltered[31]~63 (
	.dataa(!\A_ctrl_shift_rot~q ),
	.datab(!\A_data_ram_ld_align_sign_bit~q ),
	.datac(!\A_ctrl_ld_signed~q ),
	.datad(!\A_slow_inst_sel~q ),
	.datae(!\A_shift_rot_result[31]~q ),
	.dataf(!\A_slow_inst_result[31]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[31]~63_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[31]~63 .extended_lut = "off";
defparam \A_wr_data_unfiltered[31]~63 .lut_mask = 64'h7FBFFFFFFFFFFFFF;
defparam \A_wr_data_unfiltered[31]~63 .shared_arith = "off";

cyclonev_lcell_comb \A_wr_data_unfiltered[31]~64 (
	.dataa(!\A_ctrl_mul_lsw~q ),
	.datab(!\A_inst_result[31]~q ),
	.datac(!\A_wr_data_unfiltered[29]~32_combout ),
	.datad(!\A_mul_result[31]~q ),
	.datae(!\A_wr_data_unfiltered[31]~63_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_wr_data_unfiltered[31]~64_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_wr_data_unfiltered[31]~64 .extended_lut = "off";
defparam \A_wr_data_unfiltered[31]~64 .lut_mask = 64'h7BFFFFFF7BFFFFFF;
defparam \A_wr_data_unfiltered[31]~64 .shared_arith = "off";

dffeas \W_wr_data[31] (
	.clk(clk_clk),
	.d(\A_wr_data_unfiltered[31]~64_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\W_wr_data[31]~q ),
	.prn(vcc));
defparam \W_wr_data[31] .is_wysiwyg = "true";
defparam \W_wr_data[31] .power_up = "low";

cyclonev_lcell_comb \D_src1_reg[31]~15 (
	.dataa(!\embedded_system_nios2_qsys_0_register_bank_a|the_altsyncram|auto_generated|q_b[31] ),
	.datab(!\W_wr_data[31]~q ),
	.datac(!\M_alu_result[31]~q ),
	.datad(!\A_wr_data_unfiltered[31]~64_combout ),
	.datae(!\E_src1[7]~0_combout ),
	.dataf(!\E_src1[7]~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src1_reg[31]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src1_reg[31]~15 .extended_lut = "off";
defparam \D_src1_reg[31]~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \D_src1_reg[31]~15 .shared_arith = "off";

dffeas \E_src1[31] (
	.clk(clk_clk),
	.d(\D_src1_reg[31]~15_combout ),
	.asdata(\E_alu_result[31]~combout ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\Equal296~0_combout ),
	.sload(\D_src1_hazard_E~combout ),
	.ena(\A_stall~combout ),
	.q(\E_src1[31]~q ),
	.prn(vcc));
defparam \E_src1[31] .is_wysiwyg = "true";
defparam \E_src1[31] .power_up = "low";

cyclonev_lcell_comb \Add17~37 (
	.dataa(!\E_ctrl_alu_signed_comparison~q ),
	.datab(!\E_ctrl_alu_subtract~q ),
	.datac(gnd),
	.datad(!\E_src2[31]~q ),
	.datae(gnd),
	.dataf(!\E_src1[31]~q ),
	.datag(gnd),
	.cin(\Add17~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~37_sumout ),
	.cout(\Add17~38 ),
	.shareout());
defparam \Add17~37 .extended_lut = "off";
defparam \Add17~37 .lut_mask = 64'h000055AA00009966;
defparam \Add17~37 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~61 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add17~37_sumout ),
	.datac(!\D_src2_reg[0]~28_combout ),
	.datad(!\E_alu_result~30_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~61_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~61 .extended_lut = "off";
defparam \D_src2_reg[31]~61 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \D_src2_reg[31]~61 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~62 (
	.dataa(!\D_src2_reg[5]~3_combout ),
	.datab(!\D_src2_reg[5]~4_combout ),
	.datac(!\D_src2_reg[13]~8_combout ),
	.datad(!\W_wr_data[31]~q ),
	.datae(!\A_wr_data_unfiltered[31]~64_combout ),
	.dataf(!\M_alu_result[31]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~62_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~62 .extended_lut = "off";
defparam \D_src2_reg[31]~62 .lut_mask = 64'h6FFFFFFFFFFFFFFF;
defparam \D_src2_reg[31]~62 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[31]~6 (
	.dataa(!\D_iw[21]~q ),
	.datab(!\D_ctrl_unsigned_lo_imm16~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[31]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[31]~6 .extended_lut = "off";
defparam \D_src2[31]~6 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \D_src2[31]~6 .shared_arith = "off";

cyclonev_lcell_comb \D_src2[31]~7 (
	.dataa(!\D_ctrl_src2_choose_imm~q ),
	.datab(!\D_src2_reg[0]~55_combout ),
	.datac(!\D_src2_reg[31]~61_combout ),
	.datad(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.datae(!\D_src2_reg[31]~62_combout ),
	.dataf(!\D_src2[31]~6_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2[31]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2[31]~7 .extended_lut = "off";
defparam \D_src2[31]~7 .lut_mask = 64'h27FFFFFFFFFFFFFF;
defparam \D_src2[31]~7 .shared_arith = "off";

dffeas \E_src2[31] (
	.clk(clk_clk),
	.d(\D_src2[31]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2[31]~q ),
	.prn(vcc));
defparam \E_src2[31] .is_wysiwyg = "true";
defparam \E_src2[31] .power_up = "low";

cyclonev_lcell_comb \Add17~61 (
	.dataa(gnd),
	.datab(!\E_ctrl_alu_subtract~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add17~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add17~61_sumout ),
	.cout(),
	.shareout());
defparam \Add17~61 .extended_lut = "off";
defparam \Add17~61 .lut_mask = 64'h0000000000003333;
defparam \Add17~61 .shared_arith = "off";

cyclonev_lcell_comb \E_br_result~2 (
	.dataa(!\Add17~61_sumout ),
	.datab(!\E_br_result~0_combout ),
	.datac(!\E_br_result~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_br_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_br_result~2 .extended_lut = "off";
defparam \E_br_result~2 .lut_mask = 64'h2727272727272727;
defparam \E_br_result~2 .shared_arith = "off";

dffeas E_ctrl_br_cond(
	.clk(clk_clk),
	.d(\E_ctrl_br_cond_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_br_cond~q ),
	.prn(vcc));
defparam E_ctrl_br_cond.is_wysiwyg = "true";
defparam E_ctrl_br_cond.power_up = "low";

cyclonev_lcell_comb \D_ctrl_flush_pipe_always~0 (
	.dataa(!\D_iw[11]~q ),
	.datab(!\D_iw[12]~q ),
	.datac(!\D_iw[13]~q ),
	.datad(!\D_iw[14]~q ),
	.datae(!\D_iw[15]~q ),
	.dataf(!\D_iw[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_flush_pipe_always~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_flush_pipe_always~0 .extended_lut = "off";
defparam \D_ctrl_flush_pipe_always~0 .lut_mask = 64'h6996966996696996;
defparam \D_ctrl_flush_pipe_always~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_flush_pipe_always~1 (
	.dataa(!\Equal171~0_combout ),
	.datab(!\D_ctrl_flush_pipe_always~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_flush_pipe_always~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_flush_pipe_always~1 .extended_lut = "off";
defparam \D_ctrl_flush_pipe_always~1 .lut_mask = 64'h7777777777777777;
defparam \D_ctrl_flush_pipe_always~1 .shared_arith = "off";

dffeas E_ctrl_flush_pipe_always(
	.clk(clk_clk),
	.d(\D_ctrl_flush_pipe_always~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_flush_pipe_always~q ),
	.prn(vcc));
defparam E_ctrl_flush_pipe_always.is_wysiwyg = "true";
defparam E_ctrl_flush_pipe_always.power_up = "low";

cyclonev_lcell_comb \M_pipe_flush_nxt~0 (
	.dataa(!\E_valid~0_combout ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_bht_data[1]~q ),
	.datad(!\E_br_result~2_combout ),
	.datae(!\E_ctrl_br_cond~q ),
	.dataf(!\E_ctrl_flush_pipe_always~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_pipe_flush_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_pipe_flush_nxt~0 .extended_lut = "off";
defparam \M_pipe_flush_nxt~0 .lut_mask = 64'hFFFFFFFFFFFFEFFE;
defparam \M_pipe_flush_nxt~0 .shared_arith = "off";

dffeas M_pipe_flush(
	.clk(clk_clk),
	.d(\M_pipe_flush_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_pipe_flush~q ),
	.prn(vcc));
defparam M_pipe_flush.is_wysiwyg = "true";
defparam M_pipe_flush.power_up = "low";

dffeas E_wr_dst_reg_from_D(
	.clk(clk_clk),
	.d(\D_wr_dst_reg~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_wr_dst_reg_from_D~q ),
	.prn(vcc));
defparam E_wr_dst_reg_from_D.is_wysiwyg = "true";
defparam E_wr_dst_reg_from_D.power_up = "low";

cyclonev_lcell_comb \E_wr_dst_reg~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\E_hbreak_req~combout ),
	.datac(!\E_wr_dst_reg_from_D~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_wr_dst_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_wr_dst_reg~0 .extended_lut = "off";
defparam \E_wr_dst_reg~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \E_wr_dst_reg~0 .shared_arith = "off";

cyclonev_lcell_comb \E_regnum_b_cmp_F~0 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[22] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[23] ),
	.datac(!\E_dst_regnum[0]~q ),
	.datad(!\E_dst_regnum[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_b_cmp_F~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_b_cmp_F~0 .extended_lut = "off";
defparam \E_regnum_b_cmp_F~0 .lut_mask = 64'h6996699669966996;
defparam \E_regnum_b_cmp_F~0 .shared_arith = "off";

cyclonev_lcell_comb \E_regnum_b_cmp_F~1 (
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[25] ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[26] ),
	.datac(!\E_dst_regnum[3]~q ),
	.datad(!\E_dst_regnum[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_b_cmp_F~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_regnum_b_cmp_F~1 .extended_lut = "off";
defparam \E_regnum_b_cmp_F~1 .lut_mask = 64'h6996699669966996;
defparam \E_regnum_b_cmp_F~1 .shared_arith = "off";

cyclonev_lcell_comb E_regnum_b_cmp_F(
	.dataa(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[24] ),
	.datab(!\E_dst_regnum[2]~q ),
	.datac(!\E_wr_dst_reg~0_combout ),
	.datad(!\E_regnum_b_cmp_F~0_combout ),
	.datae(!\E_regnum_b_cmp_F~1_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_regnum_b_cmp_F~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam E_regnum_b_cmp_F.extended_lut = "off";
defparam E_regnum_b_cmp_F.lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam E_regnum_b_cmp_F.shared_arith = "off";

dffeas M_regnum_b_cmp_D(
	.clk(clk_clk),
	.d(\E_regnum_b_cmp_F~combout ),
	.asdata(\E_regnum_b_cmp_D~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\F_stall~combout ),
	.ena(\A_stall~combout ),
	.q(\M_regnum_b_cmp_D~q ),
	.prn(vcc));
defparam M_regnum_b_cmp_D.is_wysiwyg = "true";
defparam M_regnum_b_cmp_D.power_up = "low";

cyclonev_lcell_comb \D_data_depend~1 (
	.dataa(!\D_ctrl_a_not_src~q ),
	.datab(!\D_ctrl_b_is_dst~q ),
	.datac(!\M_ctrl_late_result~q ),
	.datad(!\M_regnum_b_cmp_D~q ),
	.datae(!\M_regnum_a_cmp_D~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_data_depend~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_data_depend~1 .extended_lut = "off";
defparam \D_data_depend~1 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \D_data_depend~1 .shared_arith = "off";

cyclonev_lcell_comb \D_dep_stall~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_issue~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_dep_stall~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_dep_stall~0 .extended_lut = "off";
defparam \D_dep_stall~0 .lut_mask = 64'h7777777777777777;
defparam \D_dep_stall~0 .shared_arith = "off";

cyclonev_lcell_comb F_stall(
	.dataa(!\A_stall~combout ),
	.datab(!\D_data_depend~0_combout ),
	.datac(!\D_data_depend~1_combout ),
	.datad(!\D_dep_stall~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_stall~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_stall.extended_lut = "off";
defparam F_stall.lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam F_stall.shared_arith = "off";

dffeas \D_iw[5] (
	.clk(clk_clk),
	.d(\F_iw[5]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[5]~q ),
	.prn(vcc));
defparam \D_iw[5] .is_wysiwyg = "true";
defparam \D_iw[5] .power_up = "low";

dffeas \E_iw[5] (
	.clk(clk_clk),
	.d(\D_iw[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_iw[5]~q ),
	.prn(vcc));
defparam \E_iw[5] .is_wysiwyg = "true";
defparam \E_iw[5] .power_up = "low";

cyclonev_lcell_comb \E_ld_st_dcache_management_bus~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[1]~q ),
	.datad(!\E_iw[4]~q ),
	.datae(!\E_iw[2]~q ),
	.dataf(!\Add17~37_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ld_st_dcache_management_bus~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ld_st_dcache_management_bus~0 .extended_lut = "off";
defparam \E_ld_st_dcache_management_bus~0 .lut_mask = 64'h5FFF3FFFFFFFFFFF;
defparam \E_ld_st_dcache_management_bus~0 .shared_arith = "off";

dffeas M_ctrl_ld_st_bypass_or_dcache_management(
	.clk(clk_clk),
	.d(\E_ld_st_dcache_management_bus~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_st_bypass_or_dcache_management~q ),
	.prn(vcc));
defparam M_ctrl_ld_st_bypass_or_dcache_management.is_wysiwyg = "true";
defparam M_ctrl_ld_st_bypass_or_dcache_management.power_up = "low";

cyclonev_lcell_comb \A_mem_stall_nxt~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_ld_st_bypass_or_dcache_management~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~0 .extended_lut = "off";
defparam \A_mem_stall_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \A_mem_stall_nxt~0 .shared_arith = "off";

dffeas M_sel_data_master(
	.clk(clk_clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_sel_data_master~q ),
	.prn(vcc));
defparam M_sel_data_master.is_wysiwyg = "true";
defparam M_sel_data_master.power_up = "low";

cyclonev_lcell_comb \M_ctrl_st_nxt~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[1]~q ),
	.datac(!\E_iw[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_ctrl_st_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_ctrl_st_nxt~0 .extended_lut = "off";
defparam \M_ctrl_st_nxt~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \M_ctrl_st_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \E_st_cache~0 (
	.dataa(!\E_iw[5]~q ),
	.datab(!\Add17~37_sumout ),
	.datac(!\M_ctrl_st_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_cache~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_cache~0 .extended_lut = "off";
defparam \E_st_cache~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \E_st_cache~0 .shared_arith = "off";

dffeas M_ctrl_st_non_bypass(
	.clk(clk_clk),
	.d(\E_st_cache~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_st_non_bypass~q ),
	.prn(vcc));
defparam M_ctrl_st_non_bypass.is_wysiwyg = "true";
defparam M_ctrl_st_non_bypass.power_up = "low";

cyclonev_lcell_comb \M_dc_valid_st_cache_hit~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_sel_data_master~q ),
	.datac(!\M_ctrl_st_non_bypass~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_valid_st_cache_hit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_valid_st_cache_hit~0 .extended_lut = "off";
defparam \M_dc_valid_st_cache_hit~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_dc_valid_st_cache_hit~0 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~0 (
	.dataa(!\E_valid~1_combout ),
	.datab(!\M_ctrl_mem_nxt~0_combout ),
	.datac(!\M_dc_valid_st_cache_hit~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~0 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_dc_potential_hazard_after_st_unfiltered~0 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~1 (
	.dataa(!\M_alu_result[9]~q ),
	.datab(!\M_alu_result[8]~q ),
	.datac(!\Add17~1_sumout ),
	.datad(!\Add17~5_sumout ),
	.datae(!\M_dc_potential_hazard_after_st_unfiltered~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~1 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~1 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \M_dc_potential_hazard_after_st_unfiltered~1 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~2 (
	.dataa(!\M_alu_result[6]~q ),
	.datab(!\M_alu_result[5]~q ),
	.datac(!\Add17~17_sumout ),
	.datad(!\Add17~21_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~2 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~2 .lut_mask = 64'h6996699669966996;
defparam \M_dc_potential_hazard_after_st_unfiltered~2 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~3 (
	.dataa(!\M_alu_result[4]~q ),
	.datab(!\M_alu_result[3]~q ),
	.datac(!\M_alu_result[2]~q ),
	.datad(!\Add17~25_sumout ),
	.datae(!\Add17~29_sumout ),
	.dataf(!\Add17~33_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~3 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~3 .lut_mask = 64'h6996966996696996;
defparam \M_dc_potential_hazard_after_st_unfiltered~3 .shared_arith = "off";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~4 (
	.dataa(!\M_alu_result[10]~q ),
	.datab(!\M_alu_result[7]~q ),
	.datac(!\Add17~9_sumout ),
	.datad(!\Add17~13_sumout ),
	.datae(!\M_dc_potential_hazard_after_st_unfiltered~2_combout ),
	.dataf(!\M_dc_potential_hazard_after_st_unfiltered~3_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~4 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~4 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \M_dc_potential_hazard_after_st_unfiltered~4 .shared_arith = "off";

cyclonev_lcell_comb \A_mem_stall_nxt~1 (
	.dataa(!\A_mem_stall~q ),
	.datab(!\A_mul_stall~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~1 .extended_lut = "off";
defparam \A_mem_stall_nxt~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_mem_stall_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \E_st_bus~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[1]~q ),
	.datad(!\E_iw[2]~q ),
	.datae(!\Add17~37_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_bus~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_bus~0 .extended_lut = "off";
defparam \E_st_bus~0 .lut_mask = 64'hF7FFFFFFF7FFFFFF;
defparam \E_st_bus~0 .shared_arith = "off";

dffeas M_ctrl_st_bypass(
	.clk(clk_clk),
	.d(\E_st_bus~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_st_bypass~q ),
	.prn(vcc));
defparam M_ctrl_st_bypass.is_wysiwyg = "true";
defparam M_ctrl_st_bypass.power_up = "low";

dffeas A_ctrl_st_bypass(
	.clk(clk_clk),
	.d(\M_ctrl_st_bypass~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_st_bypass~q ),
	.prn(vcc));
defparam A_ctrl_st_bypass.is_wysiwyg = "true";
defparam A_ctrl_st_bypass.power_up = "low";

cyclonev_lcell_comb \M_dc_hit~0 (
	.dataa(!\M_alu_result[11]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[3] ),
	.datac(!\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[0] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_hit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_hit~0 .extended_lut = "off";
defparam \M_dc_hit~0 .lut_mask = 64'h7B7B7B7B7B7B7B7B;
defparam \M_dc_hit~0 .shared_arith = "off";

cyclonev_lcell_comb M_dc_hit(
	.dataa(!\M_alu_result[13]~q ),
	.datab(!\M_alu_result[12]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[1] ),
	.datad(!\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[2] ),
	.datae(!\M_dc_hit~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_hit~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_dc_hit.extended_lut = "off";
defparam M_dc_hit.lut_mask = 64'h6996FFFF6996FFFF;
defparam M_dc_hit.shared_arith = "off";

cyclonev_lcell_comb \M_dc_valid_st_bypass_hit~0 (
	.dataa(!\M_ctrl_st_bypass~q ),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_dc_hit~combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_valid_st_bypass_hit~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_valid_st_bypass_hit~0 .extended_lut = "off";
defparam \M_dc_valid_st_bypass_hit~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \M_dc_valid_st_bypass_hit~0 .shared_arith = "off";

dffeas A_dc_valid_st_bypass_hit(
	.clk(clk_clk),
	.d(\M_dc_valid_st_bypass_hit~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_valid_st_bypass_hit~q ),
	.prn(vcc));
defparam A_dc_valid_st_bypass_hit.is_wysiwyg = "true";
defparam A_dc_valid_st_bypass_hit.power_up = "low";

cyclonev_lcell_comb A_st_bypass_transfer_done(
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_wr_data_cnt[3]~q ),
	.datac(!\av_wr_data_transfer~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_st_bypass_transfer_done~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_st_bypass_transfer_done.extended_lut = "off";
defparam A_st_bypass_transfer_done.lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam A_st_bypass_transfer_done.shared_arith = "off";

dffeas A_st_bypass_transfer_done_d1(
	.clk(clk_clk),
	.d(\A_st_bypass_transfer_done~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_st_bypass_transfer_done_d1~q ),
	.prn(vcc));
defparam A_st_bypass_transfer_done_d1.is_wysiwyg = "true";
defparam A_st_bypass_transfer_done_d1.power_up = "low";

dffeas A_valid(
	.clk(clk_clk),
	.d(\M_valid_from_E~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_valid~q ),
	.prn(vcc));
defparam A_valid.is_wysiwyg = "true";
defparam A_valid.power_up = "low";

cyclonev_lcell_comb \M_dc_valid_st_cache_hit~1 (
	.dataa(!\M_dc_valid_st_cache_hit~0_combout ),
	.datab(!\M_dc_hit~combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_valid_st_cache_hit~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_valid_st_cache_hit~1 .extended_lut = "off";
defparam \M_dc_valid_st_cache_hit~1 .lut_mask = 64'h7777777777777777;
defparam \M_dc_valid_st_cache_hit~1 .shared_arith = "off";

dffeas A_dc_valid_st_cache_hit(
	.clk(clk_clk),
	.d(\M_dc_valid_st_cache_hit~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_valid_st_cache_hit~q ),
	.prn(vcc));
defparam A_dc_valid_st_cache_hit.is_wysiwyg = "true";
defparam A_dc_valid_st_cache_hit.power_up = "low";

cyclonev_lcell_comb M_dc_dirty(
	.dataa(!\A_dc_valid_st_cache_hit~q ),
	.datab(!\Equal262~2_combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[4] ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_dirty~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_dc_dirty.extended_lut = "off";
defparam M_dc_dirty.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam M_dc_dirty.shared_arith = "off";

dffeas A_dc_dirty(
	.clk(clk_clk),
	.d(\M_dc_dirty~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_dirty~q ),
	.prn(vcc));
defparam A_dc_dirty.is_wysiwyg = "true";
defparam A_dc_dirty.power_up = "low";

cyclonev_lcell_comb \Equal193~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[3]~q ),
	.datad(!\E_iw[4]~q ),
	.datae(!\E_iw[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal193~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal193~0 .extended_lut = "off";
defparam \Equal193~0 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \Equal193~0 .shared_arith = "off";

dffeas M_ctrl_dc_index_wb_inv(
	.clk(clk_clk),
	.d(\Equal193~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_dc_index_wb_inv~q ),
	.prn(vcc));
defparam M_ctrl_dc_index_wb_inv.is_wysiwyg = "true";
defparam M_ctrl_dc_index_wb_inv.power_up = "low";

dffeas A_ctrl_dc_index_wb_inv(
	.clk(clk_clk),
	.d(\M_ctrl_dc_index_wb_inv~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_dc_index_wb_inv~q ),
	.prn(vcc));
defparam A_ctrl_dc_index_wb_inv.is_wysiwyg = "true";
defparam A_ctrl_dc_index_wb_inv.power_up = "low";

dffeas A_dc_hit(
	.clk(clk_clk),
	.d(\M_dc_hit~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_hit~q ),
	.prn(vcc));
defparam A_dc_hit.is_wysiwyg = "true";
defparam A_dc_hit.power_up = "low";

cyclonev_lcell_comb \E_ctrl_dc_addr_inv~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[4]~q ),
	.datad(!\E_iw[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_dc_addr_inv~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_dc_addr_inv~0 .extended_lut = "off";
defparam \E_ctrl_dc_addr_inv~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \E_ctrl_dc_addr_inv~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal181~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_ctrl_dc_addr_inv~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal181~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal181~0 .extended_lut = "off";
defparam \Equal181~0 .lut_mask = 64'h7777777777777777;
defparam \Equal181~0 .shared_arith = "off";

dffeas M_ctrl_dc_addr_wb_inv(
	.clk(clk_clk),
	.d(\Equal181~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_dc_addr_wb_inv~q ),
	.prn(vcc));
defparam M_ctrl_dc_addr_wb_inv.is_wysiwyg = "true";
defparam M_ctrl_dc_addr_wb_inv.power_up = "low";

dffeas A_ctrl_dc_addr_wb_inv(
	.clk(clk_clk),
	.d(\M_ctrl_dc_addr_wb_inv~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_dc_addr_wb_inv~q ),
	.prn(vcc));
defparam A_ctrl_dc_addr_wb_inv.is_wysiwyg = "true";
defparam A_ctrl_dc_addr_wb_inv.power_up = "low";

cyclonev_lcell_comb \Equal178~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[3]~q ),
	.datac(!\E_iw[4]~q ),
	.datad(!\E_iw[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal178~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal178~0 .extended_lut = "off";
defparam \Equal178~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \Equal178~0 .shared_arith = "off";

dffeas M_ctrl_dc_nowb_inv(
	.clk(clk_clk),
	.d(\Equal178~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_dc_nowb_inv~q ),
	.prn(vcc));
defparam M_ctrl_dc_nowb_inv.is_wysiwyg = "true";
defparam M_ctrl_dc_nowb_inv.power_up = "low";

dffeas A_ctrl_dc_nowb_inv(
	.clk(clk_clk),
	.d(\M_ctrl_dc_nowb_inv~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_dc_nowb_inv~q ),
	.prn(vcc));
defparam A_ctrl_dc_nowb_inv.is_wysiwyg = "true";
defparam A_ctrl_dc_nowb_inv.power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_offset_nxt[0]~1 (
	.dataa(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datab(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_offset_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_offset_nxt[0]~1 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_offset_nxt[0]~1 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \A_dc_xfer_rd_addr_offset_nxt[0]~1 .shared_arith = "off";

dffeas \A_dc_xfer_rd_addr_offset[0] (
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_offset_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_offset[0]~q ),
	.prn(vcc));
defparam \A_dc_xfer_rd_addr_offset[0] .is_wysiwyg = "true";
defparam \A_dc_xfer_rd_addr_offset[0] .power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_offset_nxt[1]~0 (
	.dataa(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datab(!\A_dc_xfer_rd_addr_offset[1]~q ),
	.datac(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_offset_nxt[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_offset_nxt[1]~0 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_offset_nxt[1]~0 .lut_mask = 64'hBEBEBEBEBEBEBEBE;
defparam \A_dc_xfer_rd_addr_offset_nxt[1]~0 .shared_arith = "off";

dffeas \A_dc_xfer_rd_addr_offset[1] (
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_offset_nxt[1]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_offset[1]~q ),
	.prn(vcc));
defparam \A_dc_xfer_rd_addr_offset[1] .is_wysiwyg = "true";
defparam \A_dc_xfer_rd_addr_offset[1] .power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_active_nxt~0 (
	.dataa(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datab(!\A_dc_xfer_rd_addr_done~q ),
	.datac(!\A_dc_xfer_rd_addr_active~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_active_nxt~0 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_active_nxt~0 .lut_mask = 64'hC5C5C5C5C5C5C5C5;
defparam \A_dc_xfer_rd_addr_active_nxt~0 .shared_arith = "off";

dffeas A_dc_xfer_rd_addr_active(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_active_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_active~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_addr_active.is_wysiwyg = "true";
defparam A_dc_xfer_rd_addr_active.power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_offset_nxt[2]~2 (
	.dataa(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datab(!\A_dc_xfer_rd_addr_offset[1]~q ),
	.datac(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datad(!\A_dc_xfer_rd_addr_offset[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_offset_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_offset_nxt[2]~2 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_offset_nxt[2]~2 .lut_mask = 64'hEBBEEBBEEBBEEBBE;
defparam \A_dc_xfer_rd_addr_offset_nxt[2]~2 .shared_arith = "off";

dffeas \A_dc_xfer_rd_addr_offset[2] (
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_offset_nxt[2]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_offset[2]~q ),
	.prn(vcc));
defparam \A_dc_xfer_rd_addr_offset[2] .is_wysiwyg = "true";
defparam \A_dc_xfer_rd_addr_offset[2] .power_up = "low";

cyclonev_lcell_comb A_dc_xfer_rd_addr_done_nxt(
	.dataa(!\A_dc_xfer_rd_addr_offset[1]~q ),
	.datab(!\A_dc_xfer_rd_addr_offset[0]~q ),
	.datac(!\A_dc_xfer_rd_addr_active~q ),
	.datad(!\A_dc_xfer_rd_addr_offset[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_done_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_xfer_rd_addr_done_nxt.extended_lut = "off";
defparam A_dc_xfer_rd_addr_done_nxt.lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam A_dc_xfer_rd_addr_done_nxt.shared_arith = "off";

dffeas A_dc_xfer_rd_addr_done(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_done_nxt~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_done~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_addr_done.is_wysiwyg = "true";
defparam A_dc_xfer_rd_addr_done.power_up = "low";

cyclonev_lcell_comb \A_dc_dcache_management_done_nxt~0 (
	.dataa(!\A_dc_dirty~q ),
	.datab(!\A_ctrl_dc_index_wb_inv~q ),
	.datac(!\A_dc_hit~q ),
	.datad(!\A_ctrl_dc_addr_wb_inv~q ),
	.datae(!\A_ctrl_dc_nowb_inv~q ),
	.dataf(!\A_dc_xfer_rd_addr_done~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_dcache_management_done_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_dcache_management_done_nxt~0 .extended_lut = "off";
defparam \A_dc_dcache_management_done_nxt~0 .lut_mask = 64'hFFFFFFFFFFFFFFDF;
defparam \A_dc_dcache_management_done_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb A_dc_dcache_management_done_nxt(
	.dataa(!\A_stall~combout ),
	.datab(!\A_valid~q ),
	.datac(!\A_dc_dcache_management_done_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_dcache_management_done_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_dcache_management_done_nxt.extended_lut = "off";
defparam A_dc_dcache_management_done_nxt.lut_mask = 64'hFBFBFBFBFBFBFBFB;
defparam A_dc_dcache_management_done_nxt.shared_arith = "off";

dffeas A_dc_dcache_management_done(
	.clk(clk_clk),
	.d(\A_dc_dcache_management_done_nxt~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_dcache_management_done~q ),
	.prn(vcc));
defparam A_dc_dcache_management_done.is_wysiwyg = "true";
defparam A_dc_dcache_management_done.power_up = "low";

cyclonev_lcell_comb \M_dc_potential_hazard_after_st_unfiltered~5 (
	.dataa(!\M_dc_potential_hazard_after_st_unfiltered~1_combout ),
	.datab(!\M_dc_potential_hazard_after_st_unfiltered~4_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_potential_hazard_after_st_unfiltered~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_potential_hazard_after_st_unfiltered~5 .extended_lut = "off";
defparam \M_dc_potential_hazard_after_st_unfiltered~5 .lut_mask = 64'h7777777777777777;
defparam \M_dc_potential_hazard_after_st_unfiltered~5 .shared_arith = "off";

dffeas A_dc_potential_hazard_after_st(
	.clk(clk_clk),
	.d(\M_dc_potential_hazard_after_st_unfiltered~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_potential_hazard_after_st~q ),
	.prn(vcc));
defparam A_dc_potential_hazard_after_st.is_wysiwyg = "true";
defparam A_dc_potential_hazard_after_st.power_up = "low";

cyclonev_lcell_comb \A_mem_stall_nxt~2 (
	.dataa(!\A_dc_fill_active~q ),
	.datab(!\A_dc_fill_need_extra_stall~q ),
	.datac(!\A_dc_rd_last_transfer_d1~q ),
	.datad(!\A_ld_bypass_done~combout ),
	.datae(!\A_ctrl_ld_bypass~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~2 .extended_lut = "off";
defparam \A_mem_stall_nxt~2 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \A_mem_stall_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \A_mem_stall_nxt~3 (
	.dataa(!\A_mem_stall~q ),
	.datab(!\A_dc_dcache_management_done~q ),
	.datac(!\A_dc_valid_st_cache_hit~q ),
	.datad(!\A_dc_potential_hazard_after_st~q ),
	.datae(!\A_mem_stall_nxt~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~3 .extended_lut = "off";
defparam \A_mem_stall_nxt~3 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \A_mem_stall_nxt~3 .shared_arith = "off";

cyclonev_lcell_comb \A_mem_stall_nxt~4 (
	.dataa(!\A_ctrl_st_bypass~q ),
	.datab(!\A_dc_valid_st_bypass_hit~q ),
	.datac(!\A_st_bypass_transfer_done~combout ),
	.datad(!\A_st_bypass_transfer_done_d1~q ),
	.datae(!\A_mem_stall_nxt~3_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~4 .extended_lut = "off";
defparam \A_mem_stall_nxt~4 .lut_mask = 64'hFFB8FFFFFFB8FFFF;
defparam \A_mem_stall_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \A_mem_stall_nxt~5 (
	.dataa(!\A_mem_stall_nxt~0_combout ),
	.datab(!\M_dc_potential_hazard_after_st_unfiltered~1_combout ),
	.datac(!\M_dc_potential_hazard_after_st_unfiltered~4_combout ),
	.datad(!\M_dc_want_fill~combout ),
	.datae(!\A_mem_stall_nxt~1_combout ),
	.dataf(!\A_mem_stall_nxt~4_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_stall_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_mem_stall_nxt~5 .extended_lut = "off";
defparam \A_mem_stall_nxt~5 .lut_mask = 64'h7FFFFFFFFFFFFFFF;
defparam \A_mem_stall_nxt~5 .shared_arith = "off";

dffeas A_mem_stall(
	.clk(clk_clk),
	.d(\A_mem_stall_nxt~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_mem_stall~q ),
	.prn(vcc));
defparam A_mem_stall.is_wysiwyg = "true";
defparam A_mem_stall.power_up = "low";

cyclonev_lcell_comb A_stall(
	.dataa(!\A_mem_stall~q ),
	.datab(!\A_mul_stall~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_stall~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_stall.extended_lut = "off";
defparam A_stall.lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam A_stall.shared_arith = "off";

cyclonev_lcell_comb \wait_for_one_post_bret_inst~0 (
	.dataa(!\A_stall~combout ),
	.datab(!hbreak_enabled1),
	.datac(!\E_valid~0_combout ),
	.datad(!\wait_for_one_post_bret_inst~q ),
	.datae(!\the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_single_step_mode~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wait_for_one_post_bret_inst~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wait_for_one_post_bret_inst~0 .extended_lut = "off";
defparam \wait_for_one_post_bret_inst~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \wait_for_one_post_bret_inst~0 .shared_arith = "off";

dffeas wait_for_one_post_bret_inst(
	.clk(clk_clk),
	.d(\wait_for_one_post_bret_inst~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\wait_for_one_post_bret_inst~q ),
	.prn(vcc));
defparam wait_for_one_post_bret_inst.is_wysiwyg = "true";
defparam wait_for_one_post_bret_inst.power_up = "low";

cyclonev_lcell_comb \hbreak_req~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\wait_for_one_post_bret_inst~q ),
	.datac(!\latched_oci_tb_hbreak_req~q ),
	.datad(!\the_embedded_system_nios2_qsys_0_nios2_oci|the_embedded_system_nios2_qsys_0_nios2_oci_debug|jtag_break~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_req~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_req~0 .extended_lut = "off";
defparam \hbreak_req~0 .lut_mask = 64'hEFFFEFFFEFFFEFFF;
defparam \hbreak_req~0 .shared_arith = "off";

cyclonev_lcell_comb \latched_oci_tb_hbreak_req_next~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\E_valid~0_combout ),
	.datac(!\latched_oci_tb_hbreak_req~q ),
	.datad(!\hbreak_req~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\latched_oci_tb_hbreak_req_next~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \latched_oci_tb_hbreak_req_next~0 .extended_lut = "off";
defparam \latched_oci_tb_hbreak_req_next~0 .lut_mask = 64'hA3FFA3FFA3FFA3FF;
defparam \latched_oci_tb_hbreak_req_next~0 .shared_arith = "off";

dffeas latched_oci_tb_hbreak_req(
	.clk(clk_clk),
	.d(\latched_oci_tb_hbreak_req_next~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\latched_oci_tb_hbreak_req~q ),
	.prn(vcc));
defparam latched_oci_tb_hbreak_req.is_wysiwyg = "true";
defparam latched_oci_tb_hbreak_req.power_up = "low";

cyclonev_lcell_comb \F_iw~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\latched_oci_tb_hbreak_req~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw~0 .extended_lut = "off";
defparam \F_iw~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw~0 .shared_arith = "off";

cyclonev_lcell_comb \F_iw[0]~9 (
	.dataa(!\F_iw~0_combout ),
	.datab(!\embedded_system_nios2_qsys_0_ic_data|the_altsyncram|auto_generated|q_b[0] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_iw[0]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_iw[0]~9 .extended_lut = "off";
defparam \F_iw[0]~9 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \F_iw[0]~9 .shared_arith = "off";

dffeas \D_iw[0] (
	.clk(clk_clk),
	.d(\F_iw[0]~9_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_iw[0]~q ),
	.prn(vcc));
defparam \D_iw[0] .is_wysiwyg = "true";
defparam \D_iw[0] .power_up = "low";

cyclonev_lcell_comb \Equal171~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal171~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal171~0 .extended_lut = "off";
defparam \Equal171~0 .lut_mask = 64'hFFFFFFFFBFFFFFFF;
defparam \Equal171~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_shift_rot~1 (
	.dataa(!\D_iw[14]~q ),
	.datab(!\D_iw[13]~q ),
	.datac(!\D_iw[12]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_shift_rot~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_shift_rot~1 .extended_lut = "off";
defparam \D_ctrl_shift_rot~1 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \D_ctrl_shift_rot~1 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~2 (
	.dataa(!\D_iw[16]~q ),
	.datab(!\D_iw[15]~q ),
	.datac(!\D_iw[14]~q ),
	.datad(!\D_iw[13]~q ),
	.datae(!\D_iw[12]~q ),
	.dataf(!\D_iw[11]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~2 .extended_lut = "off";
defparam \D_ctrl_late_result~2 .lut_mask = 64'hDDF5FFFFFFFFFFFF;
defparam \D_ctrl_late_result~2 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~0 (
	.dataa(!\D_iw[0]~q ),
	.datab(!\D_iw[5]~q ),
	.datac(!\D_iw[3]~q ),
	.datad(!\D_iw[1]~q ),
	.datae(!\D_iw[4]~q ),
	.dataf(!\D_iw[2]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~0 .extended_lut = "off";
defparam \D_ctrl_late_result~0 .lut_mask = 64'hFFFFF7FBFFFFFFFF;
defparam \D_ctrl_late_result~0 .shared_arith = "off";

cyclonev_lcell_comb \D_ctrl_late_result~1 (
	.dataa(!\Equal171~0_combout ),
	.datab(!\D_ctrl_shift_rot~1_combout ),
	.datac(!\D_ctrl_late_result~2_combout ),
	.datad(!\D_ctrl_late_result~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ctrl_late_result~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ctrl_late_result~1 .extended_lut = "off";
defparam \D_ctrl_late_result~1 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \D_ctrl_late_result~1 .shared_arith = "off";

dffeas E_ctrl_late_result(
	.clk(clk_clk),
	.d(\D_ctrl_late_result~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_ctrl_late_result~q ),
	.prn(vcc));
defparam E_ctrl_late_result.is_wysiwyg = "true";
defparam E_ctrl_late_result.power_up = "low";

cyclonev_lcell_comb \D_data_depend~0 (
	.dataa(!\E_ctrl_late_result~q ),
	.datab(!\D_ctrl_a_not_src~q ),
	.datac(!\E_regnum_a_cmp_D~q ),
	.datad(!\D_ctrl_b_is_dst~q ),
	.datae(!\E_regnum_b_cmp_D~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_data_depend~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_data_depend~0 .extended_lut = "off";
defparam \D_data_depend~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \D_data_depend~0 .shared_arith = "off";

cyclonev_lcell_comb D_valid(
	.dataa(!\D_data_depend~0_combout ),
	.datab(!\D_data_depend~1_combout ),
	.datac(!\D_dep_stall~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_valid~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam D_valid.extended_lut = "off";
defparam D_valid.lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam D_valid.shared_arith = "off";

dffeas E_valid_from_D(
	.clk(clk_clk),
	.d(\D_valid~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_valid_from_D~q ),
	.prn(vcc));
defparam E_valid_from_D.is_wysiwyg = "true";
defparam E_valid_from_D.power_up = "low";

cyclonev_lcell_comb \E_valid~0 (
	.dataa(!\E_valid_from_D~q ),
	.datab(!\M_pipe_flush~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid~0 .extended_lut = "off";
defparam \E_valid~0 .lut_mask = 64'h7777777777777777;
defparam \E_valid~0 .shared_arith = "off";

cyclonev_lcell_comb \E_valid~1 (
	.dataa(!\E_valid~0_combout ),
	.datab(!\E_hbreak_req~0_combout ),
	.datac(!\Equal209~0_combout ),
	.datad(!\E_hbreak_req~1_combout ),
	.datae(!\hbreak_req~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_valid~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_valid~1 .extended_lut = "off";
defparam \E_valid~1 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \E_valid~1 .shared_arith = "off";

dffeas M_valid_from_E(
	.clk(clk_clk),
	.d(\E_valid~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_valid_from_E~q ),
	.prn(vcc));
defparam M_valid_from_E.is_wysiwyg = "true";
defparam M_valid_from_E.power_up = "low";

cyclonev_lcell_comb \M_dc_want_fill~0 (
	.dataa(!\M_alu_result[13]~q ),
	.datab(!\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[2] ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_want_fill~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_want_fill~0 .extended_lut = "off";
defparam \M_dc_want_fill~0 .lut_mask = 64'h6666666666666666;
defparam \M_dc_want_fill~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ld_st_cache~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\Add17~37_sumout ),
	.datad(!\M_ctrl_ld_st_nxt~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ld_st_cache~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ld_st_cache~0 .extended_lut = "off";
defparam \E_ld_st_cache~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \E_ld_st_cache~0 .shared_arith = "off";

dffeas M_ctrl_ld_st_non_bypass(
	.clk(clk_clk),
	.d(\E_ld_st_cache~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_st_non_bypass~q ),
	.prn(vcc));
defparam M_ctrl_ld_st_non_bypass.is_wysiwyg = "true";
defparam M_ctrl_ld_st_non_bypass.power_up = "low";

cyclonev_lcell_comb \M_dc_want_fill~1 (
	.dataa(!\M_ctrl_ld_st_non_bypass~q ),
	.datab(!\M_sel_data_master~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_want_fill~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \M_dc_want_fill~1 .extended_lut = "off";
defparam \M_dc_want_fill~1 .lut_mask = 64'h7777777777777777;
defparam \M_dc_want_fill~1 .shared_arith = "off";

cyclonev_lcell_comb M_dc_want_fill(
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_alu_result[12]~q ),
	.datac(!\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[1] ),
	.datad(!\M_dc_hit~0_combout ),
	.datae(!\M_dc_want_fill~0_combout ),
	.dataf(!\M_dc_want_fill~1_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\M_dc_want_fill~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam M_dc_want_fill.extended_lut = "off";
defparam M_dc_want_fill.lut_mask = 64'hFF7DFFFFFFFFFFFF;
defparam M_dc_want_fill.shared_arith = "off";

dffeas A_dc_want_fill(
	.clk(clk_clk),
	.d(\M_dc_want_fill~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_want_fill~q ),
	.prn(vcc));
defparam A_dc_want_fill.is_wysiwyg = "true";
defparam A_dc_want_fill.power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_has_started_nxt~0 (
	.dataa(!\A_dc_xfer_rd_addr_has_started~q ),
	.datab(!\A_dc_xfer_rd_addr_starting~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_has_started_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_has_started_nxt~0 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_has_started_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \A_dc_xfer_rd_addr_has_started_nxt~0 .shared_arith = "off";

dffeas A_dc_xfer_rd_addr_has_started(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_has_started_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_addr_has_started~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_addr_has_started.is_wysiwyg = "true";
defparam A_dc_xfer_rd_addr_has_started.power_up = "low";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_starting~0 (
	.dataa(!\A_valid~q ),
	.datab(!\A_ctrl_dc_index_wb_inv~q ),
	.datac(!\A_dc_hit~q ),
	.datad(!\A_ctrl_dc_addr_wb_inv~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_starting~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_starting~0 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_starting~0 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \A_dc_xfer_rd_addr_starting~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_xfer_rd_addr_starting~1 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_dc_want_fill~q ),
	.datac(!\A_dc_dirty~q ),
	.datad(!\A_dc_xfer_rd_addr_has_started~q ),
	.datae(!\A_dc_xfer_rd_addr_starting~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_xfer_rd_addr_starting~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_xfer_rd_addr_starting~1 .extended_lut = "off";
defparam \A_dc_xfer_rd_addr_starting~1 .lut_mask = 64'hFFBFFFFFFFBFFFFF;
defparam \A_dc_xfer_rd_addr_starting~1 .shared_arith = "off";

dffeas A_dc_xfer_rd_data_starting(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_addr_starting~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_rd_data_starting~q ),
	.prn(vcc));
defparam A_dc_xfer_rd_data_starting.is_wysiwyg = "true";
defparam A_dc_xfer_rd_data_starting.power_up = "low";

dffeas A_dc_xfer_wr_starting(
	.clk(clk_clk),
	.d(\A_dc_xfer_rd_data_starting~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_xfer_wr_starting~q ),
	.prn(vcc));
defparam A_dc_xfer_wr_starting.is_wysiwyg = "true";
defparam A_dc_xfer_wr_starting.power_up = "low";

dffeas A_dc_wb_rd_addr_starting(
	.clk(clk_clk),
	.d(\A_dc_xfer_wr_starting~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_wb_rd_addr_starting~q ),
	.prn(vcc));
defparam A_dc_wb_rd_addr_starting.is_wysiwyg = "true";
defparam A_dc_wb_rd_addr_starting.power_up = "low";

dffeas A_dc_wb_rd_data_starting(
	.clk(clk_clk),
	.d(\A_dc_wb_rd_addr_starting~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_wb_rd_data_starting~q ),
	.prn(vcc));
defparam A_dc_wb_rd_data_starting.is_wysiwyg = "true";
defparam A_dc_wb_rd_data_starting.power_up = "low";

cyclonev_lcell_comb \A_dc_wb_rd_data_first_nxt~0 (
	.dataa(!d_read),
	.datab(!\A_dc_wb_rd_data_first~q ),
	.datac(!\A_dc_wb_rd_data_starting~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_rd_data_first_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_wb_rd_data_first_nxt~0 .extended_lut = "off";
defparam \A_dc_wb_rd_data_first_nxt~0 .lut_mask = 64'h4747474747474747;
defparam \A_dc_wb_rd_data_first_nxt~0 .shared_arith = "off";

dffeas A_dc_wb_rd_data_first(
	.clk(clk_clk),
	.d(\A_dc_wb_rd_data_first_nxt~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\A_dc_wb_rd_data_first~q ),
	.prn(vcc));
defparam A_dc_wb_rd_data_first.is_wysiwyg = "true";
defparam A_dc_wb_rd_data_first.power_up = "low";

cyclonev_lcell_comb \E_ld_st_bus~0 (
	.dataa(!\E_iw[0]~q ),
	.datab(!\E_iw[5]~q ),
	.datac(!\E_iw[1]~q ),
	.datad(!\E_iw[4]~q ),
	.datae(!\E_iw[2]~q ),
	.dataf(!\Add17~37_sumout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ld_st_bus~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ld_st_bus~0 .extended_lut = "off";
defparam \E_ld_st_bus~0 .lut_mask = 64'hF737FFFFFFFFFFFF;
defparam \E_ld_st_bus~0 .shared_arith = "off";

dffeas M_ctrl_ld_st_bypass(
	.clk(clk_clk),
	.d(\E_ld_st_bus~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_ld_st_bypass~q ),
	.prn(vcc));
defparam M_ctrl_ld_st_bypass.is_wysiwyg = "true";
defparam M_ctrl_ld_st_bypass.power_up = "low";

dffeas A_ctrl_ld_st_bypass(
	.clk(clk_clk),
	.d(\M_ctrl_ld_st_bypass~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ctrl_ld_st_bypass~q ),
	.prn(vcc));
defparam A_ctrl_ld_st_bypass.is_wysiwyg = "true";
defparam A_ctrl_ld_st_bypass.power_up = "low";

cyclonev_lcell_comb A_mem_bypass_pending(
	.dataa(!\A_ctrl_ld_st_bypass~q ),
	.datab(!\A_stall~combout ),
	.datac(!\A_valid~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_mem_bypass_pending~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_mem_bypass_pending.extended_lut = "off";
defparam A_mem_bypass_pending.lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam A_mem_bypass_pending.shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field[1]~0 (
	.dataa(!d_write),
	.datab(!d_read),
	.datac(!\A_dc_wb_rd_data_first~q ),
	.datad(!\A_mem_bypass_pending~combout ),
	.datae(!\A_dc_fill_starting~0_combout ),
	.dataf(!av_waitrequest),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field[1]~0 .extended_lut = "off";
defparam \d_address_offset_field[1]~0 .lut_mask = 64'hFFFFFFFFEFFFFFFF;
defparam \d_address_offset_field[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field[1]~1 (
	.dataa(!d_write),
	.datab(!d_read),
	.datac(!\A_dc_wb_rd_data_first~q ),
	.datad(!\A_mem_bypass_pending~combout ),
	.datae(!\A_dc_fill_starting~0_combout ),
	.dataf(!av_waitrequest),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field[1]~1 .extended_lut = "off";
defparam \d_address_offset_field[1]~1 .lut_mask = 64'hFFFFFFFFFFEFFFFF;
defparam \d_address_offset_field[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field_nxt[0]~0 (
	.dataa(!d_address_offset_field_0),
	.datab(!\d_address_offset_field[1]~0_combout ),
	.datac(!\d_address_offset_field[1]~1_combout ),
	.datad(!\A_mem_baddr[2]~q ),
	.datae(!\M_alu_result[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field_nxt[0]~0 .extended_lut = "off";
defparam \d_address_offset_field_nxt[0]~0 .lut_mask = 64'hBEFFFFFFBEFFFFFF;
defparam \d_address_offset_field_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field[1]~2 (
	.dataa(!\A_dc_wb_wr_starting~combout ),
	.datab(!\A_dc_wb_wr_active~q ),
	.datac(!\A_dc_fill_active~q ),
	.datad(!\A_dc_wb_active~q ),
	.datae(!\A_dc_want_fill~q ),
	.dataf(!\A_dc_fill_has_started~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field[1]~2 .extended_lut = "off";
defparam \d_address_offset_field[1]~2 .lut_mask = 64'hFFFFBFFFFFFFFFFF;
defparam \d_address_offset_field[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field[1]~3 (
	.dataa(!hold_waitrequest),
	.datab(!d_write),
	.datac(!d_read),
	.datad(!suppress_change_dest_id),
	.datae(!WideOr0),
	.dataf(!\d_address_offset_field[1]~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field[1]~3 .extended_lut = "off";
defparam \d_address_offset_field[1]~3 .lut_mask = 64'hFFFFFFFFFFFFFF7F;
defparam \d_address_offset_field[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \A_st_bypass_delayed~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\M_ctrl_st_bypass~q ),
	.datac(!\M_valid_from_E~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_st_bypass_delayed~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_st_bypass_delayed~0 .extended_lut = "off";
defparam \A_st_bypass_delayed~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \A_st_bypass_delayed~0 .shared_arith = "off";

dffeas A_st_bypass_delayed(
	.clk(clk_clk),
	.d(\A_st_bypass_delayed~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_bypass_delayed~q ),
	.prn(vcc));
defparam A_st_bypass_delayed.is_wysiwyg = "true";
defparam A_st_bypass_delayed.power_up = "low";

cyclonev_lcell_comb \A_st_bypass_delayed_started~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_st_bypass_delayed~q ),
	.datac(!\A_st_bypass_delayed_started~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_st_bypass_delayed_started~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_st_bypass_delayed_started~0 .extended_lut = "off";
defparam \A_st_bypass_delayed_started~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \A_st_bypass_delayed_started~0 .shared_arith = "off";

dffeas A_st_bypass_delayed_started(
	.clk(clk_clk),
	.d(\A_st_bypass_delayed_started~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_st_bypass_delayed_started~q ),
	.prn(vcc));
defparam A_st_bypass_delayed_started.is_wysiwyg = "true";
defparam A_st_bypass_delayed_started.power_up = "low";

cyclonev_lcell_comb \d_write_nxt~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_st_bypass_delayed~q ),
	.datac(!\A_st_bypass_delayed_started~q ),
	.datad(!\M_ctrl_st_bypass~q ),
	.datae(!\always120~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_write_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_write_nxt~0 .extended_lut = "off";
defparam \d_write_nxt~0 .lut_mask = 64'hFBFFFFFFFBFFFFFF;
defparam \d_write_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \d_write_nxt~1 (
	.dataa(!d_write),
	.datab(!\A_dc_wb_wr_starting~combout ),
	.datac(!av_waitrequest),
	.datad(!\d_write_nxt~0_combout ),
	.datae(!\A_dc_wr_data_cnt[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_write_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_write_nxt~1 .extended_lut = "off";
defparam \d_write_nxt~1 .lut_mask = 64'hFFFFF7FFFFFFF7FF;
defparam \d_write_nxt~1 .shared_arith = "off";

dffeas \A_dc_actual_tag[2] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[2] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_actual_tag[2]~q ),
	.prn(vcc));
defparam \A_dc_actual_tag[2] .is_wysiwyg = "true";
defparam \A_dc_actual_tag[2] .power_up = "low";

dffeas \A_dc_wb_tag[2] (
	.clk(clk_clk),
	.d(\A_dc_actual_tag[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_tag[2]~q ),
	.prn(vcc));
defparam \A_dc_wb_tag[2] .is_wysiwyg = "true";
defparam \A_dc_wb_tag[2] .power_up = "low";

cyclonev_lcell_comb A_dc_wb_wr_want_dmaster(
	.dataa(!\A_dc_wb_wr_starting~combout ),
	.datab(!\A_dc_wb_wr_active~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_wr_want_dmaster~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_wb_wr_want_dmaster.extended_lut = "off";
defparam A_dc_wb_wr_want_dmaster.lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam A_dc_wb_wr_want_dmaster.shared_arith = "off";

cyclonev_lcell_comb \d_address_tag_field_nxt~0 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_fill_active~q ),
	.datac(!\A_dc_fill_starting~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt~0 .extended_lut = "off";
defparam \d_address_tag_field_nxt~0 .lut_mask = 64'hFEFEFEFEFEFEFEFE;
defparam \d_address_tag_field_nxt~0 .shared_arith = "off";

dffeas \A_mem_baddr[13] (
	.clk(clk_clk),
	.d(\M_alu_result[13]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[13]~q ),
	.prn(vcc));
defparam \A_mem_baddr[13] .is_wysiwyg = "true";
defparam \A_mem_baddr[13] .power_up = "low";

cyclonev_lcell_comb \d_address_tag_field_nxt[2]~1 (
	.dataa(!\A_dc_wb_tag[2]~q ),
	.datab(!\A_dc_wb_wr_want_dmaster~combout ),
	.datac(!\d_address_tag_field_nxt~0_combout ),
	.datad(!\A_mem_baddr[13]~q ),
	.datae(!\M_alu_result[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt[2]~1 .extended_lut = "off";
defparam \d_address_tag_field_nxt[2]~1 .lut_mask = 64'h7DFFFFFF7DFFFFFF;
defparam \d_address_tag_field_nxt[2]~1 .shared_arith = "off";

dffeas \A_dc_actual_tag[1] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[1] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_actual_tag[1]~q ),
	.prn(vcc));
defparam \A_dc_actual_tag[1] .is_wysiwyg = "true";
defparam \A_dc_actual_tag[1] .power_up = "low";

dffeas \A_dc_wb_tag[1] (
	.clk(clk_clk),
	.d(\A_dc_actual_tag[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_tag[1]~q ),
	.prn(vcc));
defparam \A_dc_wb_tag[1] .is_wysiwyg = "true";
defparam \A_dc_wb_tag[1] .power_up = "low";

dffeas \A_mem_baddr[12] (
	.clk(clk_clk),
	.d(\M_alu_result[12]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[12]~q ),
	.prn(vcc));
defparam \A_mem_baddr[12] .is_wysiwyg = "true";
defparam \A_mem_baddr[12] .power_up = "low";

cyclonev_lcell_comb \d_address_tag_field_nxt[1]~2 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_tag[1]~q ),
	.datad(!\A_mem_baddr[12]~q ),
	.datae(!\M_alu_result[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt[1]~2 .extended_lut = "off";
defparam \d_address_tag_field_nxt[1]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_tag_field_nxt[1]~2 .shared_arith = "off";

dffeas \A_dc_actual_tag[0] (
	.clk(clk_clk),
	.d(\embedded_system_nios2_qsys_0_dc_tag|the_altsyncram|auto_generated|q_b[0] ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_dc_actual_tag[0]~q ),
	.prn(vcc));
defparam \A_dc_actual_tag[0] .is_wysiwyg = "true";
defparam \A_dc_actual_tag[0] .power_up = "low";

dffeas \A_dc_wb_tag[0] (
	.clk(clk_clk),
	.d(\A_dc_actual_tag[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_tag[0]~q ),
	.prn(vcc));
defparam \A_dc_wb_tag[0] .is_wysiwyg = "true";
defparam \A_dc_wb_tag[0] .power_up = "low";

dffeas \A_mem_baddr[11] (
	.clk(clk_clk),
	.d(\M_alu_result[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_baddr[11]~q ),
	.prn(vcc));
defparam \A_mem_baddr[11] .is_wysiwyg = "true";
defparam \A_mem_baddr[11] .power_up = "low";

cyclonev_lcell_comb \d_address_tag_field_nxt[0]~3 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_tag[0]~q ),
	.datad(!\A_mem_baddr[11]~q ),
	.datae(!\M_alu_result[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_tag_field_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_tag_field_nxt[0]~3 .extended_lut = "off";
defparam \d_address_tag_field_nxt[0]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_tag_field_nxt[0]~3 .shared_arith = "off";

dffeas \A_dc_wb_line[5] (
	.clk(clk_clk),
	.d(\A_mem_baddr[10]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[5]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[5] .is_wysiwyg = "true";
defparam \A_dc_wb_line[5] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[5]~0 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[5]~q ),
	.datad(!\A_mem_baddr[10]~q ),
	.datae(!\M_alu_result[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[5]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[5]~0 .extended_lut = "off";
defparam \d_address_line_field_nxt[5]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[5]~0 .shared_arith = "off";

dffeas \A_dc_wb_line[4] (
	.clk(clk_clk),
	.d(\A_mem_baddr[9]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[4]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[4] .is_wysiwyg = "true";
defparam \A_dc_wb_line[4] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[4]~1 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[4]~q ),
	.datad(!\A_mem_baddr[9]~q ),
	.datae(!\M_alu_result[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[4]~1 .extended_lut = "off";
defparam \d_address_line_field_nxt[4]~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[4]~1 .shared_arith = "off";

dffeas \A_dc_wb_line[3] (
	.clk(clk_clk),
	.d(\A_mem_baddr[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[3]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[3] .is_wysiwyg = "true";
defparam \A_dc_wb_line[3] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[3]~2 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[3]~q ),
	.datad(!\A_mem_baddr[8]~q ),
	.datae(!\M_alu_result[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[3]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[3]~2 .extended_lut = "off";
defparam \d_address_line_field_nxt[3]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[3]~2 .shared_arith = "off";

dffeas \A_dc_wb_line[2] (
	.clk(clk_clk),
	.d(\A_mem_baddr[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[2]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[2] .is_wysiwyg = "true";
defparam \A_dc_wb_line[2] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[2]~3 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[2]~q ),
	.datad(!\A_mem_baddr[7]~q ),
	.datae(!\M_alu_result[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[2]~3 .extended_lut = "off";
defparam \d_address_line_field_nxt[2]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[2]~3 .shared_arith = "off";

dffeas \A_dc_wb_line[1] (
	.clk(clk_clk),
	.d(\A_mem_baddr[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[1]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[1] .is_wysiwyg = "true";
defparam \A_dc_wb_line[1] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[1]~4 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[1]~q ),
	.datad(!\A_mem_baddr[6]~q ),
	.datae(!\M_alu_result[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[1]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[1]~4 .extended_lut = "off";
defparam \d_address_line_field_nxt[1]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[1]~4 .shared_arith = "off";

dffeas \A_dc_wb_line[0] (
	.clk(clk_clk),
	.d(\A_mem_baddr[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_xfer_rd_data_starting~q ),
	.q(\A_dc_wb_line[0]~q ),
	.prn(vcc));
defparam \A_dc_wb_line[0] .is_wysiwyg = "true";
defparam \A_dc_wb_line[0] .power_up = "low";

cyclonev_lcell_comb \d_address_line_field_nxt[0]~5 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\d_address_tag_field_nxt~0_combout ),
	.datac(!\A_dc_wb_line[0]~q ),
	.datad(!\A_mem_baddr[5]~q ),
	.datae(!\M_alu_result[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_line_field_nxt[0]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_line_field_nxt[0]~5 .extended_lut = "off";
defparam \d_address_line_field_nxt[0]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_address_line_field_nxt[0]~5 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field_nxt[2]~2 (
	.dataa(!d_address_offset_field_0),
	.datab(!d_address_offset_field_1),
	.datac(!\M_alu_result[4]~q ),
	.datad(!\d_address_offset_field[1]~0_combout ),
	.datae(!\d_address_offset_field[1]~1_combout ),
	.dataf(!\A_mem_baddr[4]~q ),
	.datag(!d_address_offset_field_2),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field_nxt[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field_nxt[2]~2 .extended_lut = "on";
defparam \d_address_offset_field_nxt[2]~2 .lut_mask = 64'h6996F9F66996F9F6;
defparam \d_address_offset_field_nxt[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \d_address_offset_field_nxt[1]~1 (
	.dataa(!d_address_offset_field_1),
	.datab(!d_address_offset_field_0),
	.datac(!\d_address_offset_field[1]~0_combout ),
	.datad(!\d_address_offset_field[1]~1_combout ),
	.datae(!\A_mem_baddr[3]~q ),
	.dataf(!\M_alu_result[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_address_offset_field_nxt[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_address_offset_field_nxt[1]~1 .extended_lut = "off";
defparam \d_address_offset_field_nxt[1]~1 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \d_address_offset_field_nxt[1]~1 .shared_arith = "off";

cyclonev_lcell_comb A_dc_wb_update_av_writedata(
	.dataa(!hold_waitrequest),
	.datab(!\A_dc_wb_wr_starting~combout ),
	.datac(!\A_dc_wb_wr_active~q ),
	.datad(!suppress_change_dest_id),
	.datae(!WideOr0),
	.dataf(!\A_dc_wr_data_cnt[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_wb_update_av_writedata~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam A_dc_wb_update_av_writedata.extended_lut = "off";
defparam A_dc_wb_update_av_writedata.lut_mask = 64'hFEFFFFFFFFFFFFFF;
defparam A_dc_wb_update_av_writedata.shared_arith = "off";

dffeas \E_src2_reg[3] (
	.clk(clk_clk),
	.d(\D_src2_reg[3]~23_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[3]~q ),
	.prn(vcc));
defparam \E_src2_reg[3] .is_wysiwyg = "true";
defparam \E_src2_reg[3] .power_up = "low";

dffeas \E_src2_reg[11] (
	.clk(clk_clk),
	.d(\D_src2_reg[11]~120_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[11]~q ),
	.prn(vcc));
defparam \E_src2_reg[11] .is_wysiwyg = "true";
defparam \E_src2_reg[11] .power_up = "low";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'h7777777777777777;
defparam \Equal0~0 .shared_arith = "off";

dffeas \M_st_data[11] (
	.clk(clk_clk),
	.d(\E_src2_reg[3]~q ),
	.asdata(\E_src2_reg[11]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[11]~q ),
	.prn(vcc));
defparam \M_st_data[11] .is_wysiwyg = "true";
defparam \M_st_data[11] .power_up = "low";

dffeas \A_st_data[11] (
	.clk(clk_clk),
	.d(\M_st_data[11]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[11]~q ),
	.prn(vcc));
defparam \A_st_data[11] .is_wysiwyg = "true";
defparam \A_st_data[11] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[11]~0 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[11] ),
	.datad(!\A_st_data[11]~q ),
	.datae(!\M_st_data[11]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[11]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[11]~0 .extended_lut = "off";
defparam \d_writedata_nxt[11]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[11]~0 .shared_arith = "off";

cyclonev_lcell_comb \d_writedata[14]~0 (
	.dataa(!hold_waitrequest),
	.datab(!\A_dc_wb_wr_starting~combout ),
	.datac(!\A_dc_wb_wr_active~q ),
	.datad(!suppress_change_dest_id),
	.datae(!WideOr0),
	.dataf(!\A_dc_wr_data_cnt[3]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata[14]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata[14]~0 .extended_lut = "off";
defparam \d_writedata[14]~0 .lut_mask = 64'hFFFFFFFFFFFFFFF7;
defparam \d_writedata[14]~0 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\Add17~53_sumout ),
	.datad(!\Add17~57_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en~0 .extended_lut = "off";
defparam \E_mem_byte_en~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \E_mem_byte_en~0 .shared_arith = "off";

dffeas \M_mem_byte_en[0] (
	.clk(clk_clk),
	.d(\E_mem_byte_en~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_mem_byte_en[0]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[0] .is_wysiwyg = "true";
defparam \M_mem_byte_en[0] .power_up = "low";

dffeas \A_mem_byte_en[0] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_byte_en[0]~q ),
	.prn(vcc));
defparam \A_mem_byte_en[0] .is_wysiwyg = "true";
defparam \A_mem_byte_en[0] .power_up = "low";

cyclonev_lcell_comb \d_byteenable_nxt[1]~0 (
	.dataa(!\A_dc_wb_wr_want_dmaster~combout ),
	.datab(!\A_dc_fill_active~q ),
	.datac(!\A_dc_fill_starting~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_byteenable_nxt[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_byteenable_nxt[1]~0 .extended_lut = "off";
defparam \d_byteenable_nxt[1]~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \d_byteenable_nxt[1]~0 .shared_arith = "off";

cyclonev_lcell_comb \d_byteenable_nxt[0]~1 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_mem_byte_en[0]~q ),
	.datac(!\M_mem_byte_en[0]~q ),
	.datad(!\d_byteenable_nxt[1]~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_byteenable_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_byteenable_nxt[0]~1 .extended_lut = "off";
defparam \d_byteenable_nxt[0]~1 .lut_mask = 64'hBF1FBF1FBF1FBF1F;
defparam \d_byteenable_nxt[0]~1 .shared_arith = "off";

dffeas \E_src2_reg[2] (
	.clk(clk_clk),
	.d(\D_src2_reg[2]~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[2]~q ),
	.prn(vcc));
defparam \E_src2_reg[2] .is_wysiwyg = "true";
defparam \E_src2_reg[2] .power_up = "low";

dffeas \E_src2_reg[10] (
	.clk(clk_clk),
	.d(\D_src2_reg[10]~116_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[10]~q ),
	.prn(vcc));
defparam \E_src2_reg[10] .is_wysiwyg = "true";
defparam \E_src2_reg[10] .power_up = "low";

dffeas \M_st_data[10] (
	.clk(clk_clk),
	.d(\E_src2_reg[2]~q ),
	.asdata(\E_src2_reg[10]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[10]~q ),
	.prn(vcc));
defparam \M_st_data[10] .is_wysiwyg = "true";
defparam \M_st_data[10] .power_up = "low";

dffeas \A_st_data[10] (
	.clk(clk_clk),
	.d(\M_st_data[10]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[10]~q ),
	.prn(vcc));
defparam \A_st_data[10] .is_wysiwyg = "true";
defparam \A_st_data[10] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[10]~1 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[10] ),
	.datad(!\A_st_data[10]~q ),
	.datae(!\M_st_data[10]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[10]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[10]~1 .extended_lut = "off";
defparam \d_writedata_nxt[10]~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[10]~1 .shared_arith = "off";

dffeas \E_src2_reg[1] (
	.clk(clk_clk),
	.d(\D_src2_reg[1]~25_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[1]~q ),
	.prn(vcc));
defparam \E_src2_reg[1] .is_wysiwyg = "true";
defparam \E_src2_reg[1] .power_up = "low";

dffeas \E_src2_reg[9] (
	.clk(clk_clk),
	.d(\D_src2_reg[9]~112_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[9]~q ),
	.prn(vcc));
defparam \E_src2_reg[9] .is_wysiwyg = "true";
defparam \E_src2_reg[9] .power_up = "low";

dffeas \M_st_data[9] (
	.clk(clk_clk),
	.d(\E_src2_reg[1]~q ),
	.asdata(\E_src2_reg[9]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[9]~q ),
	.prn(vcc));
defparam \M_st_data[9] .is_wysiwyg = "true";
defparam \M_st_data[9] .power_up = "low";

dffeas \A_st_data[9] (
	.clk(clk_clk),
	.d(\M_st_data[9]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[9]~q ),
	.prn(vcc));
defparam \A_st_data[9] .is_wysiwyg = "true";
defparam \A_st_data[9] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[9]~2 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[9] ),
	.datad(!\A_st_data[9]~q ),
	.datae(!\M_st_data[9]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[9]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[9]~2 .extended_lut = "off";
defparam \d_writedata_nxt[9]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[9]~2 .shared_arith = "off";

dffeas \E_src2_reg[0] (
	.clk(clk_clk),
	.d(\D_src2_reg[0]~27_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[0]~q ),
	.prn(vcc));
defparam \E_src2_reg[0] .is_wysiwyg = "true";
defparam \E_src2_reg[0] .power_up = "low";

dffeas \E_src2_reg[8] (
	.clk(clk_clk),
	.d(\D_src2_reg[8]~108_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[8]~q ),
	.prn(vcc));
defparam \E_src2_reg[8] .is_wysiwyg = "true";
defparam \E_src2_reg[8] .power_up = "low";

dffeas \M_st_data[8] (
	.clk(clk_clk),
	.d(\E_src2_reg[0]~q ),
	.asdata(\E_src2_reg[8]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[8]~q ),
	.prn(vcc));
defparam \M_st_data[8] .is_wysiwyg = "true";
defparam \M_st_data[8] .power_up = "low";

dffeas \A_st_data[8] (
	.clk(clk_clk),
	.d(\M_st_data[8]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[8]~q ),
	.prn(vcc));
defparam \A_st_data[8] .is_wysiwyg = "true";
defparam \A_st_data[8] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[8]~3 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[8] ),
	.datad(!\A_st_data[8]~q ),
	.datae(!\M_st_data[8]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[8]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[8]~3 .extended_lut = "off";
defparam \d_writedata_nxt[8]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[8]~3 .shared_arith = "off";

dffeas \E_src2_reg[5] (
	.clk(clk_clk),
	.d(\D_src2_reg[5]~19_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[5]~q ),
	.prn(vcc));
defparam \E_src2_reg[5] .is_wysiwyg = "true";
defparam \E_src2_reg[5] .power_up = "low";

dffeas \E_src2_reg[13] (
	.clk(clk_clk),
	.d(\D_src2_reg[13]~128_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[13]~q ),
	.prn(vcc));
defparam \E_src2_reg[13] .is_wysiwyg = "true";
defparam \E_src2_reg[13] .power_up = "low";

dffeas \M_st_data[13] (
	.clk(clk_clk),
	.d(\E_src2_reg[5]~q ),
	.asdata(\E_src2_reg[13]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[13]~q ),
	.prn(vcc));
defparam \M_st_data[13] .is_wysiwyg = "true";
defparam \M_st_data[13] .power_up = "low";

dffeas \A_st_data[13] (
	.clk(clk_clk),
	.d(\M_st_data[13]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[13]~q ),
	.prn(vcc));
defparam \A_st_data[13] .is_wysiwyg = "true";
defparam \A_st_data[13] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[13]~4 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[13] ),
	.datad(!\A_st_data[13]~q ),
	.datae(!\M_st_data[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[13]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[13]~4 .extended_lut = "off";
defparam \d_writedata_nxt[13]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[13]~4 .shared_arith = "off";

dffeas \E_src2_reg[4] (
	.clk(clk_clk),
	.d(\D_src2_reg[4]~21_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[4]~q ),
	.prn(vcc));
defparam \E_src2_reg[4] .is_wysiwyg = "true";
defparam \E_src2_reg[4] .power_up = "low";

dffeas \E_src2_reg[12] (
	.clk(clk_clk),
	.d(\D_src2_reg[12]~124_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[12]~q ),
	.prn(vcc));
defparam \E_src2_reg[12] .is_wysiwyg = "true";
defparam \E_src2_reg[12] .power_up = "low";

dffeas \M_st_data[12] (
	.clk(clk_clk),
	.d(\E_src2_reg[4]~q ),
	.asdata(\E_src2_reg[12]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[12]~q ),
	.prn(vcc));
defparam \M_st_data[12] .is_wysiwyg = "true";
defparam \M_st_data[12] .power_up = "low";

dffeas \A_st_data[12] (
	.clk(clk_clk),
	.d(\M_st_data[12]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[12]~q ),
	.prn(vcc));
defparam \A_st_data[12] .is_wysiwyg = "true";
defparam \A_st_data[12] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[12]~5 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[12] ),
	.datad(!\A_st_data[12]~q ),
	.datae(!\M_st_data[12]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[12]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[12]~5 .extended_lut = "off";
defparam \d_writedata_nxt[12]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[12]~5 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[21]~78 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~14_combout ),
	.datad(!\Add17~73_sumout ),
	.datae(!\D_src2_reg[21]~29_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[21]~78_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[21]~78 .extended_lut = "off";
defparam \D_src2_reg[21]~78 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[21]~78 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[21]~30 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[21] ),
	.dataf(!\D_src2_reg[21]~78_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[21]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[21]~30 .extended_lut = "off";
defparam \D_src2_reg[21]~30 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[21]~30 .shared_arith = "off";

dffeas \E_src2_reg[21] (
	.clk(clk_clk),
	.d(\D_src2_reg[21]~30_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[21]~q ),
	.prn(vcc));
defparam \E_src2_reg[21] .is_wysiwyg = "true";
defparam \E_src2_reg[21] .power_up = "low";

dffeas \M_st_data[21] (
	.clk(clk_clk),
	.d(\E_src2_reg[5]~q ),
	.asdata(\E_src2_reg[21]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[21]~q ),
	.prn(vcc));
defparam \M_st_data[21] .is_wysiwyg = "true";
defparam \M_st_data[21] .power_up = "low";

dffeas \A_st_data[21] (
	.clk(clk_clk),
	.d(\M_st_data[21]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[21]~q ),
	.prn(vcc));
defparam \A_st_data[21] .is_wysiwyg = "true";
defparam \A_st_data[21] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[21]~6 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[21] ),
	.datad(!\A_st_data[21]~q ),
	.datae(!\M_st_data[21]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[21]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[21]~6 .extended_lut = "off";
defparam \d_writedata_nxt[21]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[21]~6 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[20]~79 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~15_combout ),
	.datad(!\Add17~77_sumout ),
	.datae(!\D_src2_reg[20]~31_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[20]~79_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[20]~79 .extended_lut = "off";
defparam \D_src2_reg[20]~79 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[20]~79 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[20]~32 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[20] ),
	.dataf(!\D_src2_reg[20]~79_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[20]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[20]~32 .extended_lut = "off";
defparam \D_src2_reg[20]~32 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[20]~32 .shared_arith = "off";

dffeas \E_src2_reg[20] (
	.clk(clk_clk),
	.d(\D_src2_reg[20]~32_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[20]~q ),
	.prn(vcc));
defparam \E_src2_reg[20] .is_wysiwyg = "true";
defparam \E_src2_reg[20] .power_up = "low";

dffeas \M_st_data[20] (
	.clk(clk_clk),
	.d(\E_src2_reg[4]~q ),
	.asdata(\E_src2_reg[20]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[20]~q ),
	.prn(vcc));
defparam \M_st_data[20] .is_wysiwyg = "true";
defparam \M_st_data[20] .power_up = "low";

dffeas \A_st_data[20] (
	.clk(clk_clk),
	.d(\M_st_data[20]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[20]~q ),
	.prn(vcc));
defparam \A_st_data[20] .is_wysiwyg = "true";
defparam \A_st_data[20] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[20]~7 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[20] ),
	.datad(!\A_st_data[20]~q ),
	.datae(!\M_st_data[20]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[20]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[20]~7 .extended_lut = "off";
defparam \d_writedata_nxt[20]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[20]~7 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[25]~80 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~16_combout ),
	.datad(!\Add17~81_sumout ),
	.datae(!\D_src2_reg[25]~33_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~80_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~80 .extended_lut = "off";
defparam \D_src2_reg[25]~80 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[25]~80 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[25]~34 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[25] ),
	.dataf(!\D_src2_reg[25]~80_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[25]~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[25]~34 .extended_lut = "off";
defparam \D_src2_reg[25]~34 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[25]~34 .shared_arith = "off";

dffeas \E_src2_reg[25] (
	.clk(clk_clk),
	.d(\D_src2_reg[25]~34_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[25]~q ),
	.prn(vcc));
defparam \E_src2_reg[25] .is_wysiwyg = "true";
defparam \E_src2_reg[25] .power_up = "low";

cyclonev_lcell_comb \E_st_data[25]~0 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[1]~q ),
	.datad(!\E_src2_reg[9]~q ),
	.datae(!\E_src2_reg[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[25]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[25]~0 .extended_lut = "off";
defparam \E_st_data[25]~0 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[25]~0 .shared_arith = "off";

dffeas \M_st_data[25] (
	.clk(clk_clk),
	.d(\E_st_data[25]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[25]~q ),
	.prn(vcc));
defparam \M_st_data[25] .is_wysiwyg = "true";
defparam \M_st_data[25] .power_up = "low";

dffeas \A_st_data[25] (
	.clk(clk_clk),
	.d(\M_st_data[25]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[25]~q ),
	.prn(vcc));
defparam \A_st_data[25] .is_wysiwyg = "true";
defparam \A_st_data[25] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[25]~8 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[25] ),
	.datad(!\A_st_data[25]~q ),
	.datae(!\M_st_data[25]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[25]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[25]~8 .extended_lut = "off";
defparam \d_writedata_nxt[25]~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[25]~8 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[17]~36 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_src2_reg[17]~35_combout ),
	.datad(!\E_alu_result[17]~combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[17] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[17]~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[17]~36 .extended_lut = "off";
defparam \D_src2_reg[17]~36 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[17]~36 .shared_arith = "off";

dffeas \E_src2_reg[17] (
	.clk(clk_clk),
	.d(\D_src2_reg[17]~36_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[17]~q ),
	.prn(vcc));
defparam \E_src2_reg[17] .is_wysiwyg = "true";
defparam \E_src2_reg[17] .power_up = "low";

dffeas \M_st_data[17] (
	.clk(clk_clk),
	.d(\E_src2_reg[1]~q ),
	.asdata(\E_src2_reg[17]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[17]~q ),
	.prn(vcc));
defparam \M_st_data[17] .is_wysiwyg = "true";
defparam \M_st_data[17] .power_up = "low";

dffeas \A_st_data[17] (
	.clk(clk_clk),
	.d(\M_st_data[17]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[17]~q ),
	.prn(vcc));
defparam \A_st_data[17] .is_wysiwyg = "true";
defparam \A_st_data[17] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[17]~9 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[17] ),
	.datad(!\A_st_data[17]~q ),
	.datae(!\M_st_data[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[17]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[17]~9 .extended_lut = "off";
defparam \d_writedata_nxt[17]~9 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[17]~9 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[24]~81 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~18_combout ),
	.datad(!\Add17~89_sumout ),
	.datae(!\D_src2_reg[24]~37_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~81_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~81 .extended_lut = "off";
defparam \D_src2_reg[24]~81 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[24]~81 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[24]~38 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[24] ),
	.dataf(!\D_src2_reg[24]~81_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[24]~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[24]~38 .extended_lut = "off";
defparam \D_src2_reg[24]~38 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[24]~38 .shared_arith = "off";

dffeas \E_src2_reg[24] (
	.clk(clk_clk),
	.d(\D_src2_reg[24]~38_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[24]~q ),
	.prn(vcc));
defparam \E_src2_reg[24] .is_wysiwyg = "true";
defparam \E_src2_reg[24] .power_up = "low";

cyclonev_lcell_comb \E_st_data[24]~1 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[0]~q ),
	.datad(!\E_src2_reg[8]~q ),
	.datae(!\E_src2_reg[24]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[24]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[24]~1 .extended_lut = "off";
defparam \E_st_data[24]~1 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[24]~1 .shared_arith = "off";

dffeas \M_st_data[24] (
	.clk(clk_clk),
	.d(\E_st_data[24]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[24]~q ),
	.prn(vcc));
defparam \M_st_data[24] .is_wysiwyg = "true";
defparam \M_st_data[24] .power_up = "low";

dffeas \A_st_data[24] (
	.clk(clk_clk),
	.d(\M_st_data[24]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[24]~q ),
	.prn(vcc));
defparam \A_st_data[24] .is_wysiwyg = "true";
defparam \A_st_data[24] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[24]~10 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[24] ),
	.datad(!\A_st_data[24]~q ),
	.datae(!\M_st_data[24]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[24]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[24]~10 .extended_lut = "off";
defparam \d_writedata_nxt[24]~10 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[24]~10 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[16]~40 (
	.dataa(!\D_src2_reg[5]~1_combout ),
	.datab(!\D_src2_reg[5]~2_combout ),
	.datac(!\D_src2_reg[16]~39_combout ),
	.datad(!\E_alu_result[16]~combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[16] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[16]~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[16]~40 .extended_lut = "off";
defparam \D_src2_reg[16]~40 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \D_src2_reg[16]~40 .shared_arith = "off";

dffeas \E_src2_reg[16] (
	.clk(clk_clk),
	.d(\D_src2_reg[16]~40_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[16]~q ),
	.prn(vcc));
defparam \E_src2_reg[16] .is_wysiwyg = "true";
defparam \E_src2_reg[16] .power_up = "low";

dffeas \M_st_data[16] (
	.clk(clk_clk),
	.d(\E_src2_reg[0]~q ),
	.asdata(\E_src2_reg[16]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[16]~q ),
	.prn(vcc));
defparam \M_st_data[16] .is_wysiwyg = "true";
defparam \M_st_data[16] .power_up = "low";

dffeas \A_st_data[16] (
	.clk(clk_clk),
	.d(\M_st_data[16]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[16]~q ),
	.prn(vcc));
defparam \A_st_data[16] .is_wysiwyg = "true";
defparam \A_st_data[16] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[16]~11 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[16] ),
	.datad(!\A_st_data[16]~q ),
	.datae(!\M_st_data[16]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[16]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[16]~11 .extended_lut = "off";
defparam \d_writedata_nxt[16]~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[16]~11 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~82 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~20_combout ),
	.datad(!\Add17~97_sumout ),
	.datae(!\D_src2_reg[27]~41_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~82_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~82 .extended_lut = "off";
defparam \D_src2_reg[27]~82 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[27]~82 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[27]~42 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[27] ),
	.dataf(!\D_src2_reg[27]~82_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[27]~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[27]~42 .extended_lut = "off";
defparam \D_src2_reg[27]~42 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[27]~42 .shared_arith = "off";

dffeas \E_src2_reg[27] (
	.clk(clk_clk),
	.d(\D_src2_reg[27]~42_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[27]~q ),
	.prn(vcc));
defparam \E_src2_reg[27] .is_wysiwyg = "true";
defparam \E_src2_reg[27] .power_up = "low";

cyclonev_lcell_comb \E_st_data[27]~2 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[3]~q ),
	.datad(!\E_src2_reg[11]~q ),
	.datae(!\E_src2_reg[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[27]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[27]~2 .extended_lut = "off";
defparam \E_st_data[27]~2 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[27]~2 .shared_arith = "off";

dffeas \M_st_data[27] (
	.clk(clk_clk),
	.d(\E_st_data[27]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[27]~q ),
	.prn(vcc));
defparam \M_st_data[27] .is_wysiwyg = "true";
defparam \M_st_data[27] .power_up = "low";

dffeas \A_st_data[27] (
	.clk(clk_clk),
	.d(\M_st_data[27]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[27]~q ),
	.prn(vcc));
defparam \A_st_data[27] .is_wysiwyg = "true";
defparam \A_st_data[27] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[27]~12 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[27] ),
	.datad(!\A_st_data[27]~q ),
	.datae(!\M_st_data[27]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[27]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[27]~12 .extended_lut = "off";
defparam \d_writedata_nxt[27]~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[27]~12 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[19]~83 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~21_combout ),
	.datad(!\Add17~101_sumout ),
	.datae(!\D_src2_reg[19]~43_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[19]~83_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[19]~83 .extended_lut = "off";
defparam \D_src2_reg[19]~83 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[19]~83 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[19]~44 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[19] ),
	.dataf(!\D_src2_reg[19]~83_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[19]~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[19]~44 .extended_lut = "off";
defparam \D_src2_reg[19]~44 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[19]~44 .shared_arith = "off";

dffeas \E_src2_reg[19] (
	.clk(clk_clk),
	.d(\D_src2_reg[19]~44_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[19]~q ),
	.prn(vcc));
defparam \E_src2_reg[19] .is_wysiwyg = "true";
defparam \E_src2_reg[19] .power_up = "low";

dffeas \M_st_data[19] (
	.clk(clk_clk),
	.d(\E_src2_reg[3]~q ),
	.asdata(\E_src2_reg[19]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[19]~q ),
	.prn(vcc));
defparam \M_st_data[19] .is_wysiwyg = "true";
defparam \M_st_data[19] .power_up = "low";

dffeas \A_st_data[19] (
	.clk(clk_clk),
	.d(\M_st_data[19]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[19]~q ),
	.prn(vcc));
defparam \A_st_data[19] .is_wysiwyg = "true";
defparam \A_st_data[19] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[19]~13 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[19] ),
	.datad(!\A_st_data[19]~q ),
	.datae(!\M_st_data[19]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[19]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[19]~13 .extended_lut = "off";
defparam \d_writedata_nxt[19]~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[19]~13 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[26]~84 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~22_combout ),
	.datad(!\Add17~105_sumout ),
	.datae(!\D_src2_reg[26]~45_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~84_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~84 .extended_lut = "off";
defparam \D_src2_reg[26]~84 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[26]~84 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[26]~46 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[26] ),
	.dataf(!\D_src2_reg[26]~84_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[26]~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[26]~46 .extended_lut = "off";
defparam \D_src2_reg[26]~46 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[26]~46 .shared_arith = "off";

dffeas \E_src2_reg[26] (
	.clk(clk_clk),
	.d(\D_src2_reg[26]~46_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[26]~q ),
	.prn(vcc));
defparam \E_src2_reg[26] .is_wysiwyg = "true";
defparam \E_src2_reg[26] .power_up = "low";

cyclonev_lcell_comb \E_st_data[26]~3 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[2]~q ),
	.datad(!\E_src2_reg[10]~q ),
	.datae(!\E_src2_reg[26]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[26]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[26]~3 .extended_lut = "off";
defparam \E_st_data[26]~3 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[26]~3 .shared_arith = "off";

dffeas \M_st_data[26] (
	.clk(clk_clk),
	.d(\E_st_data[26]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[26]~q ),
	.prn(vcc));
defparam \M_st_data[26] .is_wysiwyg = "true";
defparam \M_st_data[26] .power_up = "low";

dffeas \A_st_data[26] (
	.clk(clk_clk),
	.d(\M_st_data[26]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[26]~q ),
	.prn(vcc));
defparam \A_st_data[26] .is_wysiwyg = "true";
defparam \A_st_data[26] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[26]~14 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[26] ),
	.datad(!\A_st_data[26]~q ),
	.datae(!\M_st_data[26]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[26]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[26]~14 .extended_lut = "off";
defparam \d_writedata_nxt[26]~14 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[26]~14 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[18]~85 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~23_combout ),
	.datad(!\Add17~109_sumout ),
	.datae(!\D_src2_reg[18]~47_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[18]~85_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[18]~85 .extended_lut = "off";
defparam \D_src2_reg[18]~85 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[18]~85 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[18]~48 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[18] ),
	.dataf(!\D_src2_reg[18]~85_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[18]~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[18]~48 .extended_lut = "off";
defparam \D_src2_reg[18]~48 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[18]~48 .shared_arith = "off";

dffeas \E_src2_reg[18] (
	.clk(clk_clk),
	.d(\D_src2_reg[18]~48_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[18]~q ),
	.prn(vcc));
defparam \E_src2_reg[18] .is_wysiwyg = "true";
defparam \E_src2_reg[18] .power_up = "low";

dffeas \M_st_data[18] (
	.clk(clk_clk),
	.d(\E_src2_reg[2]~q ),
	.asdata(\E_src2_reg[18]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[18]~q ),
	.prn(vcc));
defparam \M_st_data[18] .is_wysiwyg = "true";
defparam \M_st_data[18] .power_up = "low";

dffeas \A_st_data[18] (
	.clk(clk_clk),
	.d(\M_st_data[18]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[18]~q ),
	.prn(vcc));
defparam \A_st_data[18] .is_wysiwyg = "true";
defparam \A_st_data[18] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[18]~15 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[18] ),
	.datad(!\A_st_data[18]~q ),
	.datae(!\M_st_data[18]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[18]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[18]~15 .extended_lut = "off";
defparam \d_writedata_nxt[18]~15 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[18]~15 .shared_arith = "off";

dffeas \E_src2_reg[7] (
	.clk(clk_clk),
	.d(\D_src2_reg[7]~15_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[7]~q ),
	.prn(vcc));
defparam \E_src2_reg[7] .is_wysiwyg = "true";
defparam \E_src2_reg[7] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[23]~86 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~24_combout ),
	.datad(!\Add17~113_sumout ),
	.datae(!\D_src2_reg[23]~49_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~86_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~86 .extended_lut = "off";
defparam \D_src2_reg[23]~86 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[23]~86 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[23]~50 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[23] ),
	.dataf(!\D_src2_reg[23]~86_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[23]~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[23]~50 .extended_lut = "off";
defparam \D_src2_reg[23]~50 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[23]~50 .shared_arith = "off";

dffeas \E_src2_reg[23] (
	.clk(clk_clk),
	.d(\D_src2_reg[23]~50_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[23]~q ),
	.prn(vcc));
defparam \E_src2_reg[23] .is_wysiwyg = "true";
defparam \E_src2_reg[23] .power_up = "low";

dffeas \M_st_data[23] (
	.clk(clk_clk),
	.d(\E_src2_reg[7]~q ),
	.asdata(\E_src2_reg[23]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[23]~q ),
	.prn(vcc));
defparam \M_st_data[23] .is_wysiwyg = "true";
defparam \M_st_data[23] .power_up = "low";

dffeas \A_st_data[23] (
	.clk(clk_clk),
	.d(\M_st_data[23]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[23]~q ),
	.prn(vcc));
defparam \A_st_data[23] .is_wysiwyg = "true";
defparam \A_st_data[23] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[23]~16 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[23] ),
	.datad(!\A_st_data[23]~q ),
	.datae(!\M_st_data[23]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[23]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[23]~16 .extended_lut = "off";
defparam \d_writedata_nxt[23]~16 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[23]~16 .shared_arith = "off";

dffeas \E_src2_reg[15] (
	.clk(clk_clk),
	.d(\D_src2_reg[15]~104_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[15]~q ),
	.prn(vcc));
defparam \E_src2_reg[15] .is_wysiwyg = "true";
defparam \E_src2_reg[15] .power_up = "low";

dffeas \M_st_data[15] (
	.clk(clk_clk),
	.d(\E_src2_reg[7]~q ),
	.asdata(\E_src2_reg[15]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[15]~q ),
	.prn(vcc));
defparam \M_st_data[15] .is_wysiwyg = "true";
defparam \M_st_data[15] .power_up = "low";

dffeas \A_st_data[15] (
	.clk(clk_clk),
	.d(\M_st_data[15]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[15]~q ),
	.prn(vcc));
defparam \A_st_data[15] .is_wysiwyg = "true";
defparam \A_st_data[15] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[15]~17 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[15] ),
	.datad(!\A_st_data[15]~q ),
	.datae(!\M_st_data[15]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[15]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[15]~17 .extended_lut = "off";
defparam \d_writedata_nxt[15]~17 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[15]~17 .shared_arith = "off";

dffeas \E_src2_reg[6] (
	.clk(clk_clk),
	.d(\D_src2_reg[6]~17_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[6]~q ),
	.prn(vcc));
defparam \E_src2_reg[6] .is_wysiwyg = "true";
defparam \E_src2_reg[6] .power_up = "low";

cyclonev_lcell_comb \D_src2_reg[22]~87 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~26_combout ),
	.datad(!\Add17~121_sumout ),
	.datae(!\D_src2_reg[22]~52_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[22]~87_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[22]~87 .extended_lut = "off";
defparam \D_src2_reg[22]~87 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[22]~87 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[22]~53 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[22] ),
	.dataf(!\D_src2_reg[22]~87_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[22]~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[22]~53 .extended_lut = "off";
defparam \D_src2_reg[22]~53 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[22]~53 .shared_arith = "off";

dffeas \E_src2_reg[22] (
	.clk(clk_clk),
	.d(\D_src2_reg[22]~53_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[22]~q ),
	.prn(vcc));
defparam \E_src2_reg[22] .is_wysiwyg = "true";
defparam \E_src2_reg[22] .power_up = "low";

dffeas \M_st_data[22] (
	.clk(clk_clk),
	.d(\E_src2_reg[6]~q ),
	.asdata(\E_src2_reg[22]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\E_iw[4]~q ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[22]~q ),
	.prn(vcc));
defparam \M_st_data[22] .is_wysiwyg = "true";
defparam \M_st_data[22] .power_up = "low";

dffeas \A_st_data[22] (
	.clk(clk_clk),
	.d(\M_st_data[22]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[22]~q ),
	.prn(vcc));
defparam \A_st_data[22] .is_wysiwyg = "true";
defparam \A_st_data[22] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[22]~18 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[22] ),
	.datad(!\A_st_data[22]~q ),
	.datae(!\M_st_data[22]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[22]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[22]~18 .extended_lut = "off";
defparam \d_writedata_nxt[22]~18 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[22]~18 .shared_arith = "off";

dffeas \E_src2_reg[14] (
	.clk(clk_clk),
	.d(\D_src2_reg[14]~100_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[14]~q ),
	.prn(vcc));
defparam \E_src2_reg[14] .is_wysiwyg = "true";
defparam \E_src2_reg[14] .power_up = "low";

dffeas \M_st_data[14] (
	.clk(clk_clk),
	.d(\E_src2_reg[6]~q ),
	.asdata(\E_src2_reg[14]~q ),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\Equal0~0_combout ),
	.ena(\A_stall~combout ),
	.q(\M_st_data[14]~q ),
	.prn(vcc));
defparam \M_st_data[14] .is_wysiwyg = "true";
defparam \M_st_data[14] .power_up = "low";

dffeas \A_st_data[14] (
	.clk(clk_clk),
	.d(\M_st_data[14]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[14]~q ),
	.prn(vcc));
defparam \A_st_data[14] .is_wysiwyg = "true";
defparam \A_st_data[14] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[14]~19 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[14] ),
	.datad(!\A_st_data[14]~q ),
	.datae(!\M_st_data[14]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[14]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[14]~19 .extended_lut = "off";
defparam \d_writedata_nxt[14]~19 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[14]~19 .shared_arith = "off";

cyclonev_lcell_comb \A_ld_bypass_delayed~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\M_valid_from_E~q ),
	.datac(!\M_ctrl_ld_bypass~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_ld_bypass_delayed~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_ld_bypass_delayed~0 .extended_lut = "off";
defparam \A_ld_bypass_delayed~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \A_ld_bypass_delayed~0 .shared_arith = "off";

dffeas A_ld_bypass_delayed(
	.clk(clk_clk),
	.d(\A_ld_bypass_delayed~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_ld_bypass_delayed~q ),
	.prn(vcc));
defparam A_ld_bypass_delayed.is_wysiwyg = "true";
defparam A_ld_bypass_delayed.power_up = "low";

cyclonev_lcell_comb \A_ld_bypass_delayed_started~0 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\A_ld_bypass_delayed~q ),
	.datac(!\A_ld_bypass_delayed_started~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_ld_bypass_delayed_started~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_ld_bypass_delayed_started~0 .extended_lut = "off";
defparam \A_ld_bypass_delayed_started~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \A_ld_bypass_delayed_started~0 .shared_arith = "off";

dffeas A_ld_bypass_delayed_started(
	.clk(clk_clk),
	.d(\A_ld_bypass_delayed_started~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(\A_stall~combout ),
	.sload(gnd),
	.ena(vcc),
	.q(\A_ld_bypass_delayed_started~q ),
	.prn(vcc));
defparam A_ld_bypass_delayed_started.is_wysiwyg = "true";
defparam A_ld_bypass_delayed_started.power_up = "low";

cyclonev_lcell_comb \d_read_nxt~0 (
	.dataa(!\A_dc_want_fill~q ),
	.datab(!\A_dc_fill_has_started~q ),
	.datac(!\A_ld_bypass_delayed~q ),
	.datad(!\A_ld_bypass_delayed_started~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_read_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_read_nxt~0 .extended_lut = "off";
defparam \d_read_nxt~0 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \d_read_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \d_read_nxt~1 (
	.dataa(!\A_dc_wb_active~q ),
	.datab(!\always120~0_combout ),
	.datac(!\M_ctrl_ld_bypass~q ),
	.datad(!\d_read_nxt~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_read_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_read_nxt~1 .extended_lut = "off";
defparam \d_read_nxt~1 .lut_mask = 64'hBFFFBFFFBFFFBFFF;
defparam \d_read_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_rd_addr_cnt_nxt[0]~3 (
	.dataa(!d_read),
	.datab(!\A_dc_fill_starting~0_combout ),
	.datac(!av_waitrequest),
	.datad(!\A_dc_rd_addr_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_addr_cnt_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_addr_cnt_nxt[0]~3 .extended_lut = "off";
defparam \A_dc_rd_addr_cnt_nxt[0]~3 .lut_mask = 64'hFF7BFF7BFF7BFF7B;
defparam \A_dc_rd_addr_cnt_nxt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_rd_addr_cnt[1]~0 (
	.dataa(!hold_waitrequest),
	.datab(!d_read),
	.datac(!\A_dc_fill_active~q ),
	.datad(!\A_dc_fill_starting~0_combout ),
	.datae(!suppress_change_dest_id),
	.dataf(!WideOr0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_addr_cnt[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_addr_cnt[1]~0 .extended_lut = "off";
defparam \A_dc_rd_addr_cnt[1]~0 .lut_mask = 64'hFFFFFFFFFFFFF7FF;
defparam \A_dc_rd_addr_cnt[1]~0 .shared_arith = "off";

dffeas \A_dc_rd_addr_cnt[0] (
	.clk(clk_clk),
	.d(\A_dc_rd_addr_cnt_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_addr_cnt[1]~0_combout ),
	.q(\A_dc_rd_addr_cnt[0]~q ),
	.prn(vcc));
defparam \A_dc_rd_addr_cnt[0] .is_wysiwyg = "true";
defparam \A_dc_rd_addr_cnt[0] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_addr_cnt_nxt[1]~2 (
	.dataa(!d_read),
	.datab(!av_waitrequest),
	.datac(!\A_dc_rd_addr_cnt[1]~q ),
	.datad(!\A_dc_rd_addr_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_addr_cnt_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_addr_cnt_nxt[1]~2 .extended_lut = "off";
defparam \A_dc_rd_addr_cnt_nxt[1]~2 .lut_mask = 64'h7FF77FF77FF77FF7;
defparam \A_dc_rd_addr_cnt_nxt[1]~2 .shared_arith = "off";

dffeas \A_dc_rd_addr_cnt[1] (
	.clk(clk_clk),
	.d(\A_dc_rd_addr_cnt_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_addr_cnt[1]~0_combout ),
	.q(\A_dc_rd_addr_cnt[1]~q ),
	.prn(vcc));
defparam \A_dc_rd_addr_cnt[1] .is_wysiwyg = "true";
defparam \A_dc_rd_addr_cnt[1] .power_up = "low";

cyclonev_lcell_comb \A_dc_rd_addr_cnt_nxt[2]~1 (
	.dataa(!d_read),
	.datab(!av_waitrequest),
	.datac(!\A_dc_rd_addr_cnt[2]~q ),
	.datad(!\A_dc_rd_addr_cnt[1]~q ),
	.datae(!\A_dc_rd_addr_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_addr_cnt_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_addr_cnt_nxt[2]~1 .extended_lut = "off";
defparam \A_dc_rd_addr_cnt_nxt[2]~1 .lut_mask = 64'hF77F7FF7F77F7FF7;
defparam \A_dc_rd_addr_cnt_nxt[2]~1 .shared_arith = "off";

dffeas \A_dc_rd_addr_cnt[2] (
	.clk(clk_clk),
	.d(\A_dc_rd_addr_cnt_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_addr_cnt[1]~0_combout ),
	.q(\A_dc_rd_addr_cnt[2]~q ),
	.prn(vcc));
defparam \A_dc_rd_addr_cnt[2] .is_wysiwyg = "true";
defparam \A_dc_rd_addr_cnt[2] .power_up = "low";

cyclonev_lcell_comb \Add15~0 (
	.dataa(!\A_dc_rd_addr_cnt[3]~q ),
	.datab(!\A_dc_rd_addr_cnt[2]~q ),
	.datac(!\A_dc_rd_addr_cnt[1]~q ),
	.datad(!\A_dc_rd_addr_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add15~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add15~0 .extended_lut = "off";
defparam \Add15~0 .lut_mask = 64'h6996699669966996;
defparam \Add15~0 .shared_arith = "off";

cyclonev_lcell_comb \A_dc_rd_addr_cnt_nxt[3]~0 (
	.dataa(!d_read),
	.datab(!\A_dc_fill_starting~0_combout ),
	.datac(!av_waitrequest),
	.datad(!\Add15~0_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\A_dc_rd_addr_cnt_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \A_dc_rd_addr_cnt_nxt[3]~0 .extended_lut = "off";
defparam \A_dc_rd_addr_cnt_nxt[3]~0 .lut_mask = 64'hDEFFDEFFDEFFDEFF;
defparam \A_dc_rd_addr_cnt_nxt[3]~0 .shared_arith = "off";

dffeas \A_dc_rd_addr_cnt[3] (
	.clk(clk_clk),
	.d(\A_dc_rd_addr_cnt_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_dc_rd_addr_cnt[1]~0_combout ),
	.q(\A_dc_rd_addr_cnt[3]~q ),
	.prn(vcc));
defparam \A_dc_rd_addr_cnt[3] .is_wysiwyg = "true";
defparam \A_dc_rd_addr_cnt[3] .power_up = "low";

cyclonev_lcell_comb \d_read_nxt~2 (
	.dataa(!d_read),
	.datab(!av_waitrequest),
	.datac(!\d_read_nxt~1_combout ),
	.datad(!\A_dc_rd_addr_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_read_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_read_nxt~2 .extended_lut = "off";
defparam \d_read_nxt~2 .lut_mask = 64'hFFDFFFDFFFDFFFDF;
defparam \d_read_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[1]~1 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\Add17~53_sumout ),
	.datad(!\Add17~57_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[1]~1 .extended_lut = "off";
defparam \E_mem_byte_en[1]~1 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \E_mem_byte_en[1]~1 .shared_arith = "off";

dffeas \M_mem_byte_en[1] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_mem_byte_en[1]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[1] .is_wysiwyg = "true";
defparam \M_mem_byte_en[1] .power_up = "low";

dffeas \A_mem_byte_en[1] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_byte_en[1]~q ),
	.prn(vcc));
defparam \A_mem_byte_en[1] .is_wysiwyg = "true";
defparam \A_mem_byte_en[1] .power_up = "low";

cyclonev_lcell_comb \d_byteenable_nxt[1]~2 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\d_byteenable_nxt[1]~0_combout ),
	.datac(!\A_mem_byte_en[1]~q ),
	.datad(!\M_mem_byte_en[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_byteenable_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_byteenable_nxt[1]~2 .extended_lut = "off";
defparam \d_byteenable_nxt[1]~2 .lut_mask = 64'h8DFF8DFF8DFF8DFF;
defparam \d_byteenable_nxt[1]~2 .shared_arith = "off";

dffeas \M_st_data[2] (
	.clk(clk_clk),
	.d(\E_src2_reg[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[2]~q ),
	.prn(vcc));
defparam \M_st_data[2] .is_wysiwyg = "true";
defparam \M_st_data[2] .power_up = "low";

dffeas \A_st_data[2] (
	.clk(clk_clk),
	.d(\M_st_data[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[2]~q ),
	.prn(vcc));
defparam \A_st_data[2] .is_wysiwyg = "true";
defparam \A_st_data[2] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[2]~20 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[2] ),
	.datad(!\A_st_data[2]~q ),
	.datae(!\M_st_data[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[2]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[2]~20 .extended_lut = "off";
defparam \d_writedata_nxt[2]~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[2]~20 .shared_arith = "off";

dffeas \M_st_data[0] (
	.clk(clk_clk),
	.d(\E_src2_reg[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[0]~q ),
	.prn(vcc));
defparam \M_st_data[0] .is_wysiwyg = "true";
defparam \M_st_data[0] .power_up = "low";

dffeas \A_st_data[0] (
	.clk(clk_clk),
	.d(\M_st_data[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[0]~q ),
	.prn(vcc));
defparam \A_st_data[0] .is_wysiwyg = "true";
defparam \A_st_data[0] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[0]~21 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[0] ),
	.datad(!\A_st_data[0]~q ),
	.datae(!\M_st_data[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[0]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[0]~21 .extended_lut = "off";
defparam \d_writedata_nxt[0]~21 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[0]~21 .shared_arith = "off";

dffeas \M_st_data[3] (
	.clk(clk_clk),
	.d(\E_src2_reg[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[3]~q ),
	.prn(vcc));
defparam \M_st_data[3] .is_wysiwyg = "true";
defparam \M_st_data[3] .power_up = "low";

dffeas \A_st_data[3] (
	.clk(clk_clk),
	.d(\M_st_data[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[3]~q ),
	.prn(vcc));
defparam \A_st_data[3] .is_wysiwyg = "true";
defparam \A_st_data[3] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[3]~22 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[3] ),
	.datad(!\A_st_data[3]~q ),
	.datae(!\M_st_data[3]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[3]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[3]~22 .extended_lut = "off";
defparam \d_writedata_nxt[3]~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[3]~22 .shared_arith = "off";

dffeas \M_st_data[1] (
	.clk(clk_clk),
	.d(\E_src2_reg[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[1]~q ),
	.prn(vcc));
defparam \M_st_data[1] .is_wysiwyg = "true";
defparam \M_st_data[1] .power_up = "low";

dffeas \A_st_data[1] (
	.clk(clk_clk),
	.d(\M_st_data[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[1]~q ),
	.prn(vcc));
defparam \A_st_data[1] .is_wysiwyg = "true";
defparam \A_st_data[1] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[1]~23 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[1] ),
	.datad(!\A_st_data[1]~q ),
	.datae(!\M_st_data[1]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[1]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[1]~23 .extended_lut = "off";
defparam \d_writedata_nxt[1]~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[1]~23 .shared_arith = "off";

cyclonev_lcell_comb \hbreak_enabled~0 (
	.dataa(!hbreak_enabled1),
	.datab(!\M_ctrl_break~q ),
	.datac(!\M_iw[14]~q ),
	.datad(!\M_op_eret~2_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\hbreak_enabled~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \hbreak_enabled~0 .extended_lut = "off";
defparam \hbreak_enabled~0 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \hbreak_enabled~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~0 (
	.dataa(!ic_fill_line_5),
	.datab(!ic_fill_line_4),
	.datac(!\F_pc[8]~q ),
	.datad(!\F_pc[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~0 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~0 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~0 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~1 (
	.dataa(!ic_fill_tag_1),
	.datab(!ic_fill_tag_0),
	.datac(!\F_pc[10]~q ),
	.datad(!\F_pc[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~1 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~1 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~1 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~2 (
	.dataa(!ic_fill_line_2),
	.datab(!ic_fill_line_1),
	.datac(!\F_pc[5]~q ),
	.datad(!\F_pc[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~2 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~2 .lut_mask = 64'h6996699669966996;
defparam \F_ic_fill_same_tag_line~2 .shared_arith = "off";

cyclonev_lcell_comb \F_ic_fill_same_tag_line~3 (
	.dataa(!ic_fill_line_3),
	.datab(!ic_fill_line_0),
	.datac(!\F_pc[6]~q ),
	.datad(!\F_pc[3]~q ),
	.datae(!\F_ic_fill_same_tag_line~1_combout ),
	.dataf(!\F_ic_fill_same_tag_line~2_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \F_ic_fill_same_tag_line~3 .extended_lut = "off";
defparam \F_ic_fill_same_tag_line~3 .lut_mask = 64'h6996FFFFFFFFFFFF;
defparam \F_ic_fill_same_tag_line~3 .shared_arith = "off";

cyclonev_lcell_comb F_ic_fill_same_tag_line(
	.dataa(!ic_fill_line_6),
	.datab(!\F_pc[9]~q ),
	.datac(!\F_ic_fill_same_tag_line~0_combout ),
	.datad(!\F_ic_fill_same_tag_line~3_combout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\F_ic_fill_same_tag_line~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam F_ic_fill_same_tag_line.extended_lut = "off";
defparam F_ic_fill_same_tag_line.lut_mask = 64'h6FFF6FFF6FFF6FFF;
defparam F_ic_fill_same_tag_line.shared_arith = "off";

dffeas D_ic_fill_same_tag_line(
	.clk(clk_clk),
	.d(\F_ic_fill_same_tag_line~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!\F_stall~combout ),
	.q(\D_ic_fill_same_tag_line~q ),
	.prn(vcc));
defparam D_ic_fill_same_tag_line.is_wysiwyg = "true";
defparam D_ic_fill_same_tag_line.power_up = "low";

cyclonev_lcell_comb \E_ctrl_invalidate_i~0 (
	.dataa(!\E_iw[12]~q ),
	.datab(!\E_iw[11]~q ),
	.datac(!\E_iw[16]~q ),
	.datad(!\E_iw[15]~q ),
	.datae(!\E_iw[13]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_invalidate_i~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_invalidate_i~0 .extended_lut = "off";
defparam \E_ctrl_invalidate_i~0 .lut_mask = 64'h9669699696696996;
defparam \E_ctrl_invalidate_i~0 .shared_arith = "off";

cyclonev_lcell_comb \E_ctrl_invalidate_i~1 (
	.dataa(!\E_iw[14]~q ),
	.datab(!\Equal209~0_combout ),
	.datac(!\E_ctrl_invalidate_i~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_ctrl_invalidate_i~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_ctrl_invalidate_i~1 .extended_lut = "off";
defparam \E_ctrl_invalidate_i~1 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \E_ctrl_invalidate_i~1 .shared_arith = "off";

dffeas M_ctrl_invalidate_i(
	.clk(clk_clk),
	.d(\E_ctrl_invalidate_i~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_ctrl_invalidate_i~q ),
	.prn(vcc));
defparam M_ctrl_invalidate_i.is_wysiwyg = "true";
defparam M_ctrl_invalidate_i.power_up = "low";

cyclonev_lcell_comb \ic_tag_clr_valid_bits_nxt~0 (
	.dataa(!\M_valid_from_E~q ),
	.datab(!\M_ctrl_invalidate_i~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_clr_valid_bits_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_clr_valid_bits_nxt~0 .extended_lut = "off";
defparam \ic_tag_clr_valid_bits_nxt~0 .lut_mask = 64'h7777777777777777;
defparam \ic_tag_clr_valid_bits_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb ic_fill_prevent_refill_nxt(
	.dataa(!\ic_fill_prevent_refill~q ),
	.datab(!\D_ic_fill_starting~0_combout ),
	.datac(!\ic_tag_clr_valid_bits_nxt~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_prevent_refill_nxt~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ic_fill_prevent_refill_nxt.extended_lut = "off";
defparam ic_fill_prevent_refill_nxt.lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam ic_fill_prevent_refill_nxt.shared_arith = "off";

dffeas ic_fill_prevent_refill(
	.clk(clk_clk),
	.d(\ic_fill_prevent_refill_nxt~combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_fill_prevent_refill~q ),
	.prn(vcc));
defparam ic_fill_prevent_refill.is_wysiwyg = "true";
defparam ic_fill_prevent_refill.power_up = "low";

cyclonev_lcell_comb \D_ic_fill_starting~0 (
	.dataa(!\M_pipe_flush~q ),
	.datab(!\D_ic_fill_same_tag_line~q ),
	.datac(!\ic_fill_prevent_refill~q ),
	.datad(!\ic_fill_active~q ),
	.datae(!\D_iw_valid~q ),
	.dataf(!\D_kill~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_ic_fill_starting~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_ic_fill_starting~0 .extended_lut = "off";
defparam \D_ic_fill_starting~0 .lut_mask = 64'hFFFFFFFFFFFFFFFD;
defparam \D_ic_fill_starting~0 .shared_arith = "off";

dffeas \ic_fill_initial_offset[2] (
	.clk(clk_clk),
	.d(\D_pc[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(\ic_fill_initial_offset[2]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[2] .power_up = "low";

dffeas D_ic_fill_starting_d1(
	.clk(clk_clk),
	.d(\D_ic_fill_starting~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\D_ic_fill_starting_d1~q ),
	.prn(vcc));
defparam D_ic_fill_starting_d1.is_wysiwyg = "true";
defparam D_ic_fill_starting_d1.power_up = "low";

dffeas \ic_fill_initial_offset[0] (
	.clk(clk_clk),
	.d(\D_pc[0]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(\ic_fill_initial_offset[0]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[0] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[0]~1 (
	.dataa(!\ic_fill_initial_offset[0]~q ),
	.datab(!\D_ic_fill_starting_d1~q ),
	.datac(!\ic_fill_dp_offset[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[0]~1 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[0]~1 .lut_mask = 64'hD1D1D1D1D1D1D1D1;
defparam \ic_fill_dp_offset_nxt[0]~1 .shared_arith = "off";

dffeas i_readdatavalid_d1(
	.clk(clk_clk),
	.d(WideOr1),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\i_readdatavalid_d1~q ),
	.prn(vcc));
defparam i_readdatavalid_d1.is_wysiwyg = "true";
defparam i_readdatavalid_d1.power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_en~0 (
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\D_ic_fill_starting_d1~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_en~0 .extended_lut = "off";
defparam \ic_fill_dp_offset_en~0 .lut_mask = 64'h7777777777777777;
defparam \ic_fill_dp_offset_en~0 .shared_arith = "off";

dffeas \ic_fill_dp_offset[0] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[0]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[0]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[0] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[0] .power_up = "low";

dffeas \ic_fill_initial_offset[1] (
	.clk(clk_clk),
	.d(\D_pc[1]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\D_ic_fill_starting~0_combout ),
	.q(\ic_fill_initial_offset[1]~q ),
	.prn(vcc));
defparam \ic_fill_initial_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_initial_offset[1] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[1]~2 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset[0]~q ),
	.datac(!\ic_fill_initial_offset[1]~q ),
	.datad(!\ic_fill_dp_offset[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[1]~2 .lut_mask = 64'h9F6F9F6F9F6F9F6F;
defparam \ic_fill_dp_offset_nxt[1]~2 .shared_arith = "off";

dffeas \ic_fill_dp_offset[1] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[1]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[1] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[1] .power_up = "low";

dffeas \ic_fill_dp_offset[2] (
	.clk(clk_clk),
	.d(\ic_fill_dp_offset_nxt[2]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_dp_offset_en~0_combout ),
	.q(\ic_fill_dp_offset[2]~q ),
	.prn(vcc));
defparam \ic_fill_dp_offset[2] .is_wysiwyg = "true";
defparam \ic_fill_dp_offset[2] .power_up = "low";

cyclonev_lcell_comb \ic_fill_dp_offset_nxt[2]~0 (
	.dataa(!\D_ic_fill_starting_d1~q ),
	.datab(!\ic_fill_dp_offset[0]~q ),
	.datac(!\ic_fill_dp_offset[1]~q ),
	.datad(!\ic_fill_initial_offset[2]~q ),
	.datae(!\ic_fill_dp_offset[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_dp_offset_nxt[2]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_dp_offset_nxt[2]~0 .extended_lut = "off";
defparam \ic_fill_dp_offset_nxt[2]~0 .lut_mask = 64'h69FF96FF69FF96FF;
defparam \ic_fill_dp_offset_nxt[2]~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_active_nxt~0 (
	.dataa(!\i_readdatavalid_d1~q ),
	.datab(!\ic_fill_initial_offset[0]~q ),
	.datac(!\ic_fill_dp_offset_nxt[0]~1_combout ),
	.datad(!\ic_fill_initial_offset[1]~q ),
	.datae(!\ic_fill_dp_offset_nxt[1]~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_active_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_active_nxt~0 .extended_lut = "off";
defparam \ic_fill_active_nxt~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \ic_fill_active_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_active_nxt~1 (
	.dataa(!\ic_fill_active~q ),
	.datab(!\D_ic_fill_starting~0_combout ),
	.datac(!\ic_fill_initial_offset[2]~q ),
	.datad(!\ic_fill_dp_offset_nxt[2]~0_combout ),
	.datae(!\ic_fill_active_nxt~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_active_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_active_nxt~1 .extended_lut = "off";
defparam \ic_fill_active_nxt~1 .lut_mask = 64'hFFFF7FF7FFFF7FF7;
defparam \ic_fill_active_nxt~1 .shared_arith = "off";

dffeas ic_fill_active(
	.clk(clk_clk),
	.d(\ic_fill_active_nxt~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\ic_fill_active~q ),
	.prn(vcc));
defparam ic_fill_active.is_wysiwyg = "true";
defparam ic_fill_active.power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[0]~3 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[0]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[0]~3 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[0]~3 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \ic_fill_ap_cnt_nxt[0]~3 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_cnt[1]~0 (
	.dataa(!src0_valid),
	.datab(!Equal1),
	.datac(!suppress_change_dest_id1),
	.datad(!WideOr01),
	.datae(!WideOr02),
	.dataf(!\D_ic_fill_starting~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt[1]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt[1]~0 .extended_lut = "off";
defparam \ic_fill_ap_cnt[1]~0 .lut_mask = 64'hD1FFFFFFFFFFFFFF;
defparam \ic_fill_ap_cnt[1]~0 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[0] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[0]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[1]~0_combout ),
	.q(\ic_fill_ap_cnt[0]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[0] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[0] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[1]~2 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[1]~q ),
	.datac(!\ic_fill_ap_cnt[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[1]~2 .lut_mask = 64'h7D7D7D7D7D7D7D7D;
defparam \ic_fill_ap_cnt_nxt[1]~2 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[1] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[1]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[1]~0_combout ),
	.q(\ic_fill_ap_cnt[1]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[1] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[1] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[2]~1 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[2]~q ),
	.datac(!\ic_fill_ap_cnt[1]~q ),
	.datad(!\ic_fill_ap_cnt[0]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[2]~1 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[2]~1 .lut_mask = 64'hD77DD77DD77DD77D;
defparam \ic_fill_ap_cnt_nxt[2]~1 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[2] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[2]~1_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[1]~0_combout ),
	.q(\ic_fill_ap_cnt[2]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[2] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[2] .power_up = "low";

cyclonev_lcell_comb \ic_fill_ap_cnt_nxt[3]~0 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!\ic_fill_ap_cnt[3]~q ),
	.datac(!\ic_fill_ap_cnt[2]~q ),
	.datad(!\ic_fill_ap_cnt[1]~q ),
	.datae(!\ic_fill_ap_cnt[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_cnt_nxt[3]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_cnt_nxt[3]~0 .extended_lut = "off";
defparam \ic_fill_ap_cnt_nxt[3]~0 .lut_mask = 64'h7DD7D77D7DD7D77D;
defparam \ic_fill_ap_cnt_nxt[3]~0 .shared_arith = "off";

dffeas \ic_fill_ap_cnt[3] (
	.clk(clk_clk),
	.d(\ic_fill_ap_cnt_nxt[3]~0_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\ic_fill_ap_cnt[1]~0_combout ),
	.q(\ic_fill_ap_cnt[3]~q ),
	.prn(vcc));
defparam \ic_fill_ap_cnt[3] .is_wysiwyg = "true";
defparam \ic_fill_ap_cnt[3] .power_up = "low";

cyclonev_lcell_comb \i_read_nxt~0 (
	.dataa(!hold_waitrequest),
	.datab(!suppress_change_dest_id1),
	.datac(!\ic_fill_active~q ),
	.datad(!\ic_fill_ap_cnt[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_read_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_read_nxt~0 .extended_lut = "off";
defparam \i_read_nxt~0 .lut_mask = 64'hFDFFFDFFFDFFFDFF;
defparam \i_read_nxt~0 .shared_arith = "off";

cyclonev_lcell_comb \i_read_nxt~1 (
	.dataa(!i_read),
	.datab(!Equal1),
	.datac(!WideOr01),
	.datad(!WideOr02),
	.datae(!\i_read_nxt~0_combout ),
	.dataf(!\D_ic_fill_starting~0_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\i_read_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \i_read_nxt~1 .extended_lut = "off";
defparam \i_read_nxt~1 .lut_mask = 64'hFFFFF7D5FFFFFFFF;
defparam \i_read_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~0 (
	.dataa(!ic_fill_line_6),
	.datab(!\D_ic_fill_starting~0_combout ),
	.datac(!\D_pc[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~0 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~0 .lut_mask = 64'h4747474747474747;
defparam \ic_tag_wraddress_nxt~0 .shared_arith = "off";

dffeas \M_st_data[6] (
	.clk(clk_clk),
	.d(\E_src2_reg[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[6]~q ),
	.prn(vcc));
defparam \M_st_data[6] .is_wysiwyg = "true";
defparam \M_st_data[6] .power_up = "low";

dffeas \A_st_data[6] (
	.clk(clk_clk),
	.d(\M_st_data[6]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[6]~q ),
	.prn(vcc));
defparam \A_st_data[6] .is_wysiwyg = "true";
defparam \A_st_data[6] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[6]~24 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[6] ),
	.datad(!\A_st_data[6]~q ),
	.datae(!\M_st_data[6]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[6]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[6]~24 .extended_lut = "off";
defparam \d_writedata_nxt[6]~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[6]~24 .shared_arith = "off";

dffeas \M_st_data[4] (
	.clk(clk_clk),
	.d(\E_src2_reg[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[4]~q ),
	.prn(vcc));
defparam \M_st_data[4] .is_wysiwyg = "true";
defparam \M_st_data[4] .power_up = "low";

dffeas \A_st_data[4] (
	.clk(clk_clk),
	.d(\M_st_data[4]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[4]~q ),
	.prn(vcc));
defparam \A_st_data[4] .is_wysiwyg = "true";
defparam \A_st_data[4] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[4]~25 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[4] ),
	.datad(!\A_st_data[4]~q ),
	.datae(!\M_st_data[4]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[4]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[4]~25 .extended_lut = "off";
defparam \d_writedata_nxt[4]~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[4]~25 .shared_arith = "off";

dffeas \M_st_data[7] (
	.clk(clk_clk),
	.d(\E_src2_reg[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[7]~q ),
	.prn(vcc));
defparam \M_st_data[7] .is_wysiwyg = "true";
defparam \M_st_data[7] .power_up = "low";

dffeas \A_st_data[7] (
	.clk(clk_clk),
	.d(\M_st_data[7]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[7]~q ),
	.prn(vcc));
defparam \A_st_data[7] .is_wysiwyg = "true";
defparam \A_st_data[7] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[7]~26 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[7] ),
	.datad(!\A_st_data[7]~q ),
	.datae(!\M_st_data[7]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[7]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[7]~26 .extended_lut = "off";
defparam \d_writedata_nxt[7]~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[7]~26 .shared_arith = "off";

dffeas \M_st_data[5] (
	.clk(clk_clk),
	.d(\E_src2_reg[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[5]~q ),
	.prn(vcc));
defparam \M_st_data[5] .is_wysiwyg = "true";
defparam \M_st_data[5] .power_up = "low";

dffeas \A_st_data[5] (
	.clk(clk_clk),
	.d(\M_st_data[5]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[5]~q ),
	.prn(vcc));
defparam \A_st_data[5] .is_wysiwyg = "true";
defparam \A_st_data[5] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[5]~27 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[5] ),
	.datad(!\A_st_data[5]~q ),
	.datae(!\M_st_data[5]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[5]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[5]~27 .extended_lut = "off";
defparam \d_writedata_nxt[5]~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[5]~27 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~1 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_5),
	.datac(!\D_pc[8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~1 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~1 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[0]~0 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!ic_fill_ap_offset_0),
	.datac(!\D_pc[0]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[0]~0 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[0]~0 .lut_mask = 64'h8D8D8D8D8D8D8D8D;
defparam \ic_fill_ap_offset_nxt[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~2 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_1),
	.datac(!\D_pc[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~2 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~2 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~2 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~3 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_0),
	.datac(!\D_pc[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~3 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~3 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~3 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[2]~1 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!ic_fill_ap_offset_0),
	.datac(!ic_fill_ap_offset_2),
	.datad(!ic_fill_ap_offset_1),
	.datae(!\D_pc[2]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[2]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[2]~1 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[2]~1 .lut_mask = 64'h6996FFFF6996FFFF;
defparam \ic_fill_ap_offset_nxt[2]~1 .shared_arith = "off";

cyclonev_lcell_comb \ic_fill_ap_offset_nxt[1]~2 (
	.dataa(!nonposted_cmd_accepted),
	.datab(!ic_fill_ap_offset_0),
	.datac(!ic_fill_ap_offset_1),
	.datad(!\D_pc[1]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_fill_ap_offset_nxt[1]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_fill_ap_offset_nxt[1]~2 .extended_lut = "off";
defparam \ic_fill_ap_offset_nxt[1]~2 .lut_mask = 64'h96FF96FF96FF96FF;
defparam \ic_fill_ap_offset_nxt[1]~2 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~4 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_4),
	.datac(!\D_pc[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~4 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~4 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~4 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~5 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_3),
	.datac(!\D_pc[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~5 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~5 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~5 .shared_arith = "off";

cyclonev_lcell_comb \ic_tag_wraddress_nxt~6 (
	.dataa(!\D_ic_fill_starting~0_combout ),
	.datab(!ic_fill_line_2),
	.datac(!\D_pc[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ic_tag_wraddress_nxt~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ic_tag_wraddress_nxt~6 .extended_lut = "off";
defparam \ic_tag_wraddress_nxt~6 .lut_mask = 64'h2727272727272727;
defparam \ic_tag_wraddress_nxt~6 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[2]~2 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\Add17~53_sumout ),
	.datad(!\Add17~57_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[2]~2 .extended_lut = "off";
defparam \E_mem_byte_en[2]~2 .lut_mask = 64'hFF7FFF7FFF7FFF7F;
defparam \E_mem_byte_en[2]~2 .shared_arith = "off";

dffeas \M_mem_byte_en[2] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[2]~2_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_mem_byte_en[2]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[2] .is_wysiwyg = "true";
defparam \M_mem_byte_en[2] .power_up = "low";

dffeas \A_mem_byte_en[2] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[2]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_byte_en[2]~q ),
	.prn(vcc));
defparam \A_mem_byte_en[2] .is_wysiwyg = "true";
defparam \A_mem_byte_en[2] .power_up = "low";

cyclonev_lcell_comb \d_byteenable_nxt[2]~3 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\d_byteenable_nxt[1]~0_combout ),
	.datac(!\M_mem_byte_en[2]~q ),
	.datad(!\A_mem_byte_en[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_byteenable_nxt[2]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_byteenable_nxt[2]~3 .extended_lut = "off";
defparam \d_byteenable_nxt[2]~3 .lut_mask = 64'h8DFF8DFF8DFF8DFF;
defparam \d_byteenable_nxt[2]~3 .shared_arith = "off";

cyclonev_lcell_comb \E_mem_byte_en[3]~3 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\Add17~53_sumout ),
	.datad(!\Add17~57_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_mem_byte_en[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_mem_byte_en[3]~3 .extended_lut = "off";
defparam \E_mem_byte_en[3]~3 .lut_mask = 64'h7FFF7FFF7FFF7FFF;
defparam \E_mem_byte_en[3]~3 .shared_arith = "off";

dffeas \M_mem_byte_en[3] (
	.clk(clk_clk),
	.d(\E_mem_byte_en[3]~3_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_mem_byte_en[3]~q ),
	.prn(vcc));
defparam \M_mem_byte_en[3] .is_wysiwyg = "true";
defparam \M_mem_byte_en[3] .power_up = "low";

dffeas \A_mem_byte_en[3] (
	.clk(clk_clk),
	.d(\M_mem_byte_en[3]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_mem_byte_en[3]~q ),
	.prn(vcc));
defparam \A_mem_byte_en[3] .is_wysiwyg = "true";
defparam \A_mem_byte_en[3] .power_up = "low";

cyclonev_lcell_comb \d_byteenable_nxt[3]~4 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\d_byteenable_nxt[1]~0_combout ),
	.datac(!\M_mem_byte_en[3]~q ),
	.datad(!\A_mem_byte_en[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_byteenable_nxt[3]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_byteenable_nxt[3]~4 .extended_lut = "off";
defparam \d_byteenable_nxt[3]~4 .lut_mask = 64'h8DFF8DFF8DFF8DFF;
defparam \d_byteenable_nxt[3]~4 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~90 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add17~37_sumout ),
	.datac(!\E_alu_result~30_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~90_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~90 .extended_lut = "off";
defparam \D_src2_reg[31]~90 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \D_src2_reg[31]~90 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[31]~75 (
	.dataa(!\D_src2_reg[0]~28_combout ),
	.datab(!\D_src2_reg[31]~62_combout ),
	.datac(!\D_src2_reg[5]~1_combout ),
	.datad(!\D_src2_reg[5]~2_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[31] ),
	.dataf(!\D_src2_reg[31]~90_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[31]~75_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[31]~75 .extended_lut = "off";
defparam \D_src2_reg[31]~75 .lut_mask = 64'hFFFFFFFFF7FFFFFF;
defparam \D_src2_reg[31]~75 .shared_arith = "off";

dffeas \E_src2_reg[31] (
	.clk(clk_clk),
	.d(\D_src2_reg[31]~75_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[31]~q ),
	.prn(vcc));
defparam \E_src2_reg[31] .is_wysiwyg = "true";
defparam \E_src2_reg[31] .power_up = "low";

cyclonev_lcell_comb \E_st_data[31]~5 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[7]~q ),
	.datad(!\E_src2_reg[15]~q ),
	.datae(!\E_src2_reg[31]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[31]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[31]~5 .extended_lut = "off";
defparam \E_st_data[31]~5 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[31]~5 .shared_arith = "off";

dffeas \M_st_data[31] (
	.clk(clk_clk),
	.d(\E_st_data[31]~5_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[31]~q ),
	.prn(vcc));
defparam \M_st_data[31] .is_wysiwyg = "true";
defparam \M_st_data[31] .power_up = "low";

dffeas \A_st_data[31] (
	.clk(clk_clk),
	.d(\M_st_data[31]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[31]~q ),
	.prn(vcc));
defparam \A_st_data[31] .is_wysiwyg = "true";
defparam \A_st_data[31] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[31]~28 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[31]~q ),
	.datad(!\A_st_data[31]~q ),
	.datae(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[31] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[31]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[31]~28 .extended_lut = "off";
defparam \d_writedata_nxt[31]~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[31]~28 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~88 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~28_combout ),
	.datad(!\Add17~129_sumout ),
	.datae(!\D_src2_reg[29]~58_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~88_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~88 .extended_lut = "off";
defparam \D_src2_reg[29]~88 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[29]~88 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[29]~74 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(!\D_src2_reg[29]~88_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[29]~74_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[29]~74 .extended_lut = "off";
defparam \D_src2_reg[29]~74 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[29]~74 .shared_arith = "off";

dffeas \E_src2_reg[29] (
	.clk(clk_clk),
	.d(\D_src2_reg[29]~74_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[29]~q ),
	.prn(vcc));
defparam \E_src2_reg[29] .is_wysiwyg = "true";
defparam \E_src2_reg[29] .power_up = "low";

cyclonev_lcell_comb \E_st_data[29]~4 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[5]~q ),
	.datad(!\E_src2_reg[13]~q ),
	.datae(!\E_src2_reg[29]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[29]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[29]~4 .extended_lut = "off";
defparam \E_st_data[29]~4 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[29]~4 .shared_arith = "off";

dffeas \M_st_data[29] (
	.clk(clk_clk),
	.d(\E_st_data[29]~4_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[29]~q ),
	.prn(vcc));
defparam \M_st_data[29] .is_wysiwyg = "true";
defparam \M_st_data[29] .power_up = "low";

dffeas \A_st_data[29] (
	.clk(clk_clk),
	.d(\M_st_data[29]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[29]~q ),
	.prn(vcc));
defparam \A_st_data[29] .is_wysiwyg = "true";
defparam \A_st_data[29] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[29]~29 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[29]~q ),
	.datad(!\A_st_data[29]~q ),
	.datae(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[29] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[29]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[29]~29 .extended_lut = "off";
defparam \d_writedata_nxt[29]~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[29]~29 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[28]~91 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\D_src2_reg[0]~28_combout ),
	.datac(!\E_alu_result~31_combout ),
	.datad(!\Add17~133_sumout ),
	.datae(!\D_src2_reg[28]~64_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~91_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~91 .extended_lut = "off";
defparam \D_src2_reg[28]~91 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[28]~91 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[28]~76 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(!\D_src2_reg[28]~91_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[28]~76_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[28]~76 .extended_lut = "off";
defparam \D_src2_reg[28]~76 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[28]~76 .shared_arith = "off";

dffeas \E_src2_reg[28] (
	.clk(clk_clk),
	.d(\D_src2_reg[28]~76_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[28]~q ),
	.prn(vcc));
defparam \E_src2_reg[28] .is_wysiwyg = "true";
defparam \E_src2_reg[28] .power_up = "low";

cyclonev_lcell_comb \E_st_data[28]~6 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[4]~q ),
	.datad(!\E_src2_reg[12]~q ),
	.datae(!\E_src2_reg[28]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[28]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[28]~6 .extended_lut = "off";
defparam \E_st_data[28]~6 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[28]~6 .shared_arith = "off";

dffeas \M_st_data[28] (
	.clk(clk_clk),
	.d(\E_st_data[28]~6_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[28]~q ),
	.prn(vcc));
defparam \M_st_data[28] .is_wysiwyg = "true";
defparam \M_st_data[28] .power_up = "low";

dffeas \A_st_data[28] (
	.clk(clk_clk),
	.d(\M_st_data[28]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[28]~q ),
	.prn(vcc));
defparam \A_st_data[28] .is_wysiwyg = "true";
defparam \A_st_data[28] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[28]~30 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[28]~q ),
	.datad(!\A_st_data[28]~q ),
	.datae(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[28] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[28]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[28]~30 .extended_lut = "off";
defparam \d_writedata_nxt[28]~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[28]~30 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[30]~89 (
	.dataa(!\E_alu_result~0_combout ),
	.datab(!\Add17~65_sumout ),
	.datac(!\D_src2_reg[0]~28_combout ),
	.datad(!\E_alu_result~29_combout ),
	.datae(!\D_src2_reg[30]~60_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~89_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~89 .extended_lut = "off";
defparam \D_src2_reg[30]~89 .lut_mask = 64'hFFFFFFFDFFFFFFFD;
defparam \D_src2_reg[30]~89 .shared_arith = "off";

cyclonev_lcell_comb \D_src2_reg[30]~77 (
	.dataa(!\D_ctrl_b_is_dst~q ),
	.datab(!\E_regnum_b_cmp_D~q ),
	.datac(!\D_src2_reg[5]~0_combout ),
	.datad(!\Equal297~0_combout ),
	.datae(!\embedded_system_nios2_qsys_0_register_bank_b|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(!\D_src2_reg[30]~89_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\D_src2_reg[30]~77_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \D_src2_reg[30]~77 .extended_lut = "off";
defparam \D_src2_reg[30]~77 .lut_mask = 64'hFFFFFFFFFFDFFFFF;
defparam \D_src2_reg[30]~77 .shared_arith = "off";

dffeas \E_src2_reg[30] (
	.clk(clk_clk),
	.d(\D_src2_reg[30]~77_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\E_src2_reg[30]~q ),
	.prn(vcc));
defparam \E_src2_reg[30] .is_wysiwyg = "true";
defparam \E_src2_reg[30] .power_up = "low";

cyclonev_lcell_comb \E_st_data[30]~7 (
	.dataa(!\E_iw[3]~q ),
	.datab(!\E_iw[4]~q ),
	.datac(!\E_src2_reg[6]~q ),
	.datad(!\E_src2_reg[14]~q ),
	.datae(!\E_src2_reg[30]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\E_st_data[30]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \E_st_data[30]~7 .extended_lut = "off";
defparam \E_st_data[30]~7 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \E_st_data[30]~7 .shared_arith = "off";

dffeas \M_st_data[30] (
	.clk(clk_clk),
	.d(\E_st_data[30]~7_combout ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\M_st_data[30]~q ),
	.prn(vcc));
defparam \M_st_data[30] .is_wysiwyg = "true";
defparam \M_st_data[30] .power_up = "low";

dffeas \A_st_data[30] (
	.clk(clk_clk),
	.d(\M_st_data[30]~q ),
	.asdata(vcc),
	.clrn(!\hq3myc14108phmpo7y7qmhbp98hy0vq~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\A_stall~combout ),
	.q(\A_st_data[30]~q ),
	.prn(vcc));
defparam \A_st_data[30] .is_wysiwyg = "true";
defparam \A_st_data[30] .power_up = "low";

cyclonev_lcell_comb \d_writedata_nxt[30]~31 (
	.dataa(!\A_mem_bypass_pending~combout ),
	.datab(!\A_dc_wb_update_av_writedata~combout ),
	.datac(!\M_st_data[30]~q ),
	.datad(!\A_st_data[30]~q ),
	.datae(!\embedded_system_nios2_qsys_0_dc_victim|the_altsyncram|auto_generated|q_b[30] ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\d_writedata_nxt[30]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \d_writedata_nxt[30]~31 .extended_lut = "off";
defparam \d_writedata_nxt[30]~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \d_writedata_nxt[30]~31 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_bht_module (
	q_b_1,
	q_b_0,
	F_stall,
	M_bht_wr_en_unfiltered,
	M_bht_wr_data_unfiltered_1,
	M_bht_ptr_unfiltered_0,
	M_bht_ptr_unfiltered_1,
	M_bht_ptr_unfiltered_2,
	M_bht_ptr_unfiltered_3,
	M_bht_ptr_unfiltered_4,
	M_bht_ptr_unfiltered_5,
	M_bht_ptr_unfiltered_6,
	M_bht_ptr_unfiltered_7,
	F_bht_ptr_nxt_0,
	F_bht_ptr_nxt_1,
	F_bht_ptr_nxt_2,
	F_bht_ptr_nxt_3,
	F_bht_ptr_nxt_4,
	F_bht_ptr_nxt_5,
	F_bht_ptr_nxt_6,
	F_bht_ptr_nxt_7,
	M_br_mispredict,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_0;
input 	F_stall;
input 	M_bht_wr_en_unfiltered;
input 	M_bht_wr_data_unfiltered_1;
input 	M_bht_ptr_unfiltered_0;
input 	M_bht_ptr_unfiltered_1;
input 	M_bht_ptr_unfiltered_2;
input 	M_bht_ptr_unfiltered_3;
input 	M_bht_ptr_unfiltered_4;
input 	M_bht_ptr_unfiltered_5;
input 	M_bht_ptr_unfiltered_6;
input 	M_bht_ptr_unfiltered_7;
input 	F_bht_ptr_nxt_0;
input 	F_bht_ptr_nxt_1;
input 	F_bht_ptr_nxt_2;
input 	F_bht_ptr_nxt_3;
input 	F_bht_ptr_nxt_4;
input 	F_bht_ptr_nxt_5;
input 	F_bht_ptr_nxt_6;
input 	F_bht_ptr_nxt_7;
input 	M_br_mispredict;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_1 the_altsyncram(
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,
q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_unconnected_wire_7,q_b_unconnected_wire_6,q_b_unconnected_wire_5,q_b_unconnected_wire_4,q_b_unconnected_wire_3,q_b_unconnected_wire_2,q_b_1,q_b_0}),
	.rden_b(F_stall),
	.wren_a(M_bht_wr_en_unfiltered),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,M_bht_wr_data_unfiltered_1,M_br_mispredict}),
	.address_a({gnd,gnd,M_bht_ptr_unfiltered_7,M_bht_ptr_unfiltered_6,M_bht_ptr_unfiltered_5,M_bht_ptr_unfiltered_4,M_bht_ptr_unfiltered_3,M_bht_ptr_unfiltered_2,M_bht_ptr_unfiltered_1,M_bht_ptr_unfiltered_0}),
	.address_b({gnd,gnd,F_bht_ptr_nxt_7,F_bht_ptr_nxt_6,F_bht_ptr_nxt_5,F_bht_ptr_nxt_4,F_bht_ptr_nxt_3,F_bht_ptr_nxt_2,F_bht_ptr_nxt_1,F_bht_ptr_nxt_0}),
	.clock0(clk_clk));

endmodule

module embedded_system_altsyncram_1 (
	q_b,
	rden_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	rden_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[9:0] address_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_9fo1 auto_generated(
	.q_b({q_b[1],q_b[0]}),
	.rden_b(rden_b),
	.wren_a(wren_a),
	.data_a({data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module embedded_system_altsyncram_9fo1 (
	q_b,
	rden_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[1:0] q_b;
input 	rden_b;
input 	wren_a;
input 	[1:0] data_a;
input 	[7:0] address_a;
input 	[7:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "embedded_system_nios2_qsys_0_bht_ram.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_bht_module:embedded_system_nios2_qsys_0_bht|altsyncram:the_altsyncram|altsyncram_9fo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 2;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 8;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 255;
defparam ram_block1a1.port_b_logical_ram_depth = 256;
defparam ram_block1a1.port_b_logical_ram_width = 2;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "C40C758C6F9E56B3BBC04C1B566B8EEE5BBC11DA8A6FB53F0F552C2614CCB91D";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "embedded_system_nios2_qsys_0_bht_ram.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_bht_module:embedded_system_nios2_qsys_0_bht|altsyncram:the_altsyncram|altsyncram_9fo1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 2;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 8;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 255;
defparam ram_block1a0.port_b_logical_ram_depth = 256;
defparam ram_block1a0.port_b_logical_ram_width = 2;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "F6602B57E2A6B55EA0889FF222FAD437FECC8623AD08233175F9DD13F8D3F521";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_dc_data_module (
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_13,
	q_b_12,
	q_b_21,
	q_b_20,
	q_b_25,
	q_b_17,
	q_b_24,
	q_b_16,
	q_b_27,
	q_b_19,
	q_b_26,
	q_b_18,
	q_b_23,
	q_b_15,
	q_b_22,
	q_b_14,
	q_b_2,
	q_b_29,
	q_b_7,
	q_b_31,
	q_b_28,
	q_b_6,
	q_b_30,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_1,
	q_b_0,
	dc_data_wr_port_en,
	dc_data_wr_port_data_11,
	dc_data_wr_port_addr_0,
	dc_data_wr_port_addr_1,
	dc_data_wr_port_addr_2,
	dc_data_wr_port_addr_3,
	dc_data_wr_port_addr_4,
	dc_data_wr_port_addr_5,
	dc_data_wr_port_addr_6,
	dc_data_wr_port_addr_7,
	dc_data_wr_port_addr_8,
	dc_data_rd_port_addr_0,
	dc_data_rd_port_addr_1,
	dc_data_rd_port_addr_2,
	dc_data_rd_port_addr_3,
	dc_data_rd_port_addr_4,
	dc_data_rd_port_addr_5,
	dc_data_rd_port_addr_6,
	dc_data_rd_port_addr_7,
	dc_data_rd_port_addr_8,
	dc_data_wr_port_data_10,
	dc_data_wr_port_data_9,
	dc_data_wr_port_data_8,
	dc_data_wr_port_data_13,
	dc_data_wr_port_data_12,
	dc_data_wr_port_data_21,
	dc_data_wr_port_data_20,
	dc_data_wr_port_data_25,
	dc_data_wr_port_data_17,
	dc_data_wr_port_data_24,
	dc_data_wr_port_data_16,
	dc_data_wr_port_data_27,
	dc_data_wr_port_data_19,
	dc_data_wr_port_data_26,
	dc_data_wr_port_data_18,
	dc_data_wr_port_data_23,
	dc_data_wr_port_data_15,
	dc_data_wr_port_data_22,
	dc_data_wr_port_data_14,
	dc_data_wr_port_data_2,
	dc_data_wr_port_data_29,
	dc_data_wr_port_data_7,
	dc_data_wr_port_data_31,
	dc_data_wr_port_data_28,
	dc_data_wr_port_data_6,
	dc_data_wr_port_data_30,
	dc_data_wr_port_data_5,
	dc_data_wr_port_data_4,
	dc_data_wr_port_data_3,
	dc_data_wr_port_data_1,
	dc_data_wr_port_data_0,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_13;
output 	q_b_12;
output 	q_b_21;
output 	q_b_20;
output 	q_b_25;
output 	q_b_17;
output 	q_b_24;
output 	q_b_16;
output 	q_b_27;
output 	q_b_19;
output 	q_b_26;
output 	q_b_18;
output 	q_b_23;
output 	q_b_15;
output 	q_b_22;
output 	q_b_14;
output 	q_b_2;
output 	q_b_29;
output 	q_b_7;
output 	q_b_31;
output 	q_b_28;
output 	q_b_6;
output 	q_b_30;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_1;
output 	q_b_0;
input 	dc_data_wr_port_en;
input 	dc_data_wr_port_data_11;
input 	dc_data_wr_port_addr_0;
input 	dc_data_wr_port_addr_1;
input 	dc_data_wr_port_addr_2;
input 	dc_data_wr_port_addr_3;
input 	dc_data_wr_port_addr_4;
input 	dc_data_wr_port_addr_5;
input 	dc_data_wr_port_addr_6;
input 	dc_data_wr_port_addr_7;
input 	dc_data_wr_port_addr_8;
input 	dc_data_rd_port_addr_0;
input 	dc_data_rd_port_addr_1;
input 	dc_data_rd_port_addr_2;
input 	dc_data_rd_port_addr_3;
input 	dc_data_rd_port_addr_4;
input 	dc_data_rd_port_addr_5;
input 	dc_data_rd_port_addr_6;
input 	dc_data_rd_port_addr_7;
input 	dc_data_rd_port_addr_8;
input 	dc_data_wr_port_data_10;
input 	dc_data_wr_port_data_9;
input 	dc_data_wr_port_data_8;
input 	dc_data_wr_port_data_13;
input 	dc_data_wr_port_data_12;
input 	dc_data_wr_port_data_21;
input 	dc_data_wr_port_data_20;
input 	dc_data_wr_port_data_25;
input 	dc_data_wr_port_data_17;
input 	dc_data_wr_port_data_24;
input 	dc_data_wr_port_data_16;
input 	dc_data_wr_port_data_27;
input 	dc_data_wr_port_data_19;
input 	dc_data_wr_port_data_26;
input 	dc_data_wr_port_data_18;
input 	dc_data_wr_port_data_23;
input 	dc_data_wr_port_data_15;
input 	dc_data_wr_port_data_22;
input 	dc_data_wr_port_data_14;
input 	dc_data_wr_port_data_2;
input 	dc_data_wr_port_data_29;
input 	dc_data_wr_port_data_7;
input 	dc_data_wr_port_data_31;
input 	dc_data_wr_port_data_28;
input 	dc_data_wr_port_data_6;
input 	dc_data_wr_port_data_30;
input 	dc_data_wr_port_data_5;
input 	dc_data_wr_port_data_4;
input 	dc_data_wr_port_data_3;
input 	dc_data_wr_port_data_1;
input 	dc_data_wr_port_data_0;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_2 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(dc_data_wr_port_en),
	.data_a({dc_data_wr_port_data_31,dc_data_wr_port_data_30,dc_data_wr_port_data_29,dc_data_wr_port_data_28,dc_data_wr_port_data_27,dc_data_wr_port_data_26,dc_data_wr_port_data_25,dc_data_wr_port_data_24,dc_data_wr_port_data_23,dc_data_wr_port_data_22,dc_data_wr_port_data_21,
dc_data_wr_port_data_20,dc_data_wr_port_data_19,dc_data_wr_port_data_18,dc_data_wr_port_data_17,dc_data_wr_port_data_16,dc_data_wr_port_data_15,dc_data_wr_port_data_14,dc_data_wr_port_data_13,dc_data_wr_port_data_12,dc_data_wr_port_data_11,dc_data_wr_port_data_10,
dc_data_wr_port_data_9,dc_data_wr_port_data_8,dc_data_wr_port_data_7,dc_data_wr_port_data_6,dc_data_wr_port_data_5,dc_data_wr_port_data_4,dc_data_wr_port_data_3,dc_data_wr_port_data_2,dc_data_wr_port_data_1,dc_data_wr_port_data_0}),
	.address_a({gnd,dc_data_wr_port_addr_8,dc_data_wr_port_addr_7,dc_data_wr_port_addr_6,dc_data_wr_port_addr_5,dc_data_wr_port_addr_4,dc_data_wr_port_addr_3,dc_data_wr_port_addr_2,dc_data_wr_port_addr_1,dc_data_wr_port_addr_0}),
	.address_b({gnd,dc_data_rd_port_addr_8,dc_data_rd_port_addr_7,dc_data_rd_port_addr_6,dc_data_rd_port_addr_5,dc_data_rd_port_addr_4,dc_data_rd_port_addr_3,dc_data_rd_port_addr_2,dc_data_rd_port_addr_1,dc_data_rd_port_addr_0}),
	.clock0(clk_clk));

endmodule

module embedded_system_altsyncram_2 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[9:0] address_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_40j1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module embedded_system_altsyncram_40j1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[8:0] address_a;
input 	[8:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 9;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 511;
defparam ram_block1a11.port_a_logical_ram_depth = 512;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 9;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 511;
defparam ram_block1a11.port_b_logical_ram_depth = 512;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 9;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 511;
defparam ram_block1a10.port_a_logical_ram_depth = 512;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 9;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 511;
defparam ram_block1a10.port_b_logical_ram_depth = 512;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 9;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 511;
defparam ram_block1a9.port_a_logical_ram_depth = 512;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 9;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 511;
defparam ram_block1a9.port_b_logical_ram_depth = 512;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 9;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 511;
defparam ram_block1a8.port_a_logical_ram_depth = 512;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 9;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 511;
defparam ram_block1a8.port_b_logical_ram_depth = 512;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 9;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 511;
defparam ram_block1a13.port_a_logical_ram_depth = 512;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 9;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 511;
defparam ram_block1a13.port_b_logical_ram_depth = 512;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 9;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 511;
defparam ram_block1a12.port_a_logical_ram_depth = 512;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 9;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 511;
defparam ram_block1a12.port_b_logical_ram_depth = 512;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 9;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 511;
defparam ram_block1a21.port_a_logical_ram_depth = 512;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 9;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 511;
defparam ram_block1a21.port_b_logical_ram_depth = 512;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 9;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 511;
defparam ram_block1a20.port_a_logical_ram_depth = 512;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 9;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 511;
defparam ram_block1a20.port_b_logical_ram_depth = 512;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 9;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 511;
defparam ram_block1a25.port_a_logical_ram_depth = 512;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 9;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 511;
defparam ram_block1a25.port_b_logical_ram_depth = 512;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 9;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 511;
defparam ram_block1a17.port_a_logical_ram_depth = 512;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 9;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 511;
defparam ram_block1a17.port_b_logical_ram_depth = 512;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 9;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 511;
defparam ram_block1a24.port_a_logical_ram_depth = 512;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 9;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 511;
defparam ram_block1a24.port_b_logical_ram_depth = 512;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 9;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 511;
defparam ram_block1a16.port_a_logical_ram_depth = 512;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 9;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 511;
defparam ram_block1a16.port_b_logical_ram_depth = 512;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 9;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 511;
defparam ram_block1a27.port_a_logical_ram_depth = 512;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 9;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 511;
defparam ram_block1a27.port_b_logical_ram_depth = 512;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 9;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 511;
defparam ram_block1a19.port_a_logical_ram_depth = 512;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 9;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 511;
defparam ram_block1a19.port_b_logical_ram_depth = 512;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 9;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 511;
defparam ram_block1a26.port_a_logical_ram_depth = 512;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 9;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 511;
defparam ram_block1a26.port_b_logical_ram_depth = 512;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 9;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 511;
defparam ram_block1a18.port_a_logical_ram_depth = 512;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 9;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 511;
defparam ram_block1a18.port_b_logical_ram_depth = 512;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 9;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 511;
defparam ram_block1a23.port_a_logical_ram_depth = 512;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 9;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 511;
defparam ram_block1a23.port_b_logical_ram_depth = 512;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 9;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 511;
defparam ram_block1a15.port_a_logical_ram_depth = 512;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 9;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 511;
defparam ram_block1a15.port_b_logical_ram_depth = 512;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 9;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 511;
defparam ram_block1a22.port_a_logical_ram_depth = 512;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 9;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 511;
defparam ram_block1a22.port_b_logical_ram_depth = 512;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 9;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 511;
defparam ram_block1a14.port_a_logical_ram_depth = 512;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 9;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 511;
defparam ram_block1a14.port_b_logical_ram_depth = 512;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 9;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 511;
defparam ram_block1a2.port_a_logical_ram_depth = 512;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 9;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 511;
defparam ram_block1a2.port_b_logical_ram_depth = 512;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 9;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 511;
defparam ram_block1a29.port_a_logical_ram_depth = 512;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 9;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 511;
defparam ram_block1a29.port_b_logical_ram_depth = 512;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 9;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 511;
defparam ram_block1a7.port_a_logical_ram_depth = 512;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 9;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 511;
defparam ram_block1a7.port_b_logical_ram_depth = 512;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 9;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 511;
defparam ram_block1a31.port_a_logical_ram_depth = 512;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 9;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 511;
defparam ram_block1a31.port_b_logical_ram_depth = 512;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 9;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 511;
defparam ram_block1a28.port_a_logical_ram_depth = 512;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 9;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 511;
defparam ram_block1a28.port_b_logical_ram_depth = 512;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 9;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 511;
defparam ram_block1a6.port_a_logical_ram_depth = 512;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 9;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 511;
defparam ram_block1a6.port_b_logical_ram_depth = 512;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 9;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 511;
defparam ram_block1a30.port_a_logical_ram_depth = 512;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 9;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 511;
defparam ram_block1a30.port_b_logical_ram_depth = 512;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 9;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 511;
defparam ram_block1a5.port_a_logical_ram_depth = 512;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 9;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 511;
defparam ram_block1a5.port_b_logical_ram_depth = 512;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 9;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 511;
defparam ram_block1a4.port_a_logical_ram_depth = 512;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 9;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 511;
defparam ram_block1a4.port_b_logical_ram_depth = 512;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 9;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 511;
defparam ram_block1a3.port_a_logical_ram_depth = 512;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 9;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 511;
defparam ram_block1a3.port_b_logical_ram_depth = 512;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 9;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 511;
defparam ram_block1a1.port_a_logical_ram_depth = 512;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 9;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 511;
defparam ram_block1a1.port_b_logical_ram_depth = 512;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_data_module:embedded_system_nios2_qsys_0_dc_data|altsyncram:the_altsyncram|altsyncram_40j1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 9;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 511;
defparam ram_block1a0.port_a_logical_ram_depth = 512;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 9;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 511;
defparam ram_block1a0.port_b_logical_ram_depth = 512;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_dc_tag_module (
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_0,
	q_b_4,
	dc_tag_wr_port_en,
	dc_tag_wr_port_data_1,
	dc_tag_wr_port_addr_0,
	dc_tag_wr_port_addr_1,
	dc_tag_wr_port_addr_2,
	dc_tag_wr_port_addr_3,
	dc_tag_wr_port_addr_4,
	dc_tag_wr_port_addr_5,
	dc_tag_rd_port_addr_0,
	dc_tag_rd_port_addr_1,
	dc_tag_rd_port_addr_2,
	dc_tag_rd_port_addr_3,
	dc_tag_rd_port_addr_4,
	dc_tag_rd_port_addr_5,
	dc_tag_wr_port_data_2,
	dc_tag_wr_port_data_3,
	dc_tag_wr_port_data_0,
	dc_tag_wr_port_data_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_0;
output 	q_b_4;
input 	dc_tag_wr_port_en;
input 	dc_tag_wr_port_data_1;
input 	dc_tag_wr_port_addr_0;
input 	dc_tag_wr_port_addr_1;
input 	dc_tag_wr_port_addr_2;
input 	dc_tag_wr_port_addr_3;
input 	dc_tag_wr_port_addr_4;
input 	dc_tag_wr_port_addr_5;
input 	dc_tag_rd_port_addr_0;
input 	dc_tag_rd_port_addr_1;
input 	dc_tag_rd_port_addr_2;
input 	dc_tag_rd_port_addr_3;
input 	dc_tag_rd_port_addr_4;
input 	dc_tag_rd_port_addr_5;
input 	dc_tag_wr_port_data_2;
input 	dc_tag_wr_port_data_3;
input 	dc_tag_wr_port_data_0;
input 	dc_tag_wr_port_data_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_3 the_altsyncram(
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,
q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_unconnected_wire_7,q_b_unconnected_wire_6,q_b_unconnected_wire_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(dc_tag_wr_port_en),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dc_tag_wr_port_data_4,dc_tag_wr_port_data_3,dc_tag_wr_port_data_2,dc_tag_wr_port_data_1,dc_tag_wr_port_data_0}),
	.address_a({gnd,gnd,gnd,gnd,dc_tag_wr_port_addr_5,dc_tag_wr_port_addr_4,dc_tag_wr_port_addr_3,dc_tag_wr_port_addr_2,dc_tag_wr_port_addr_1,dc_tag_wr_port_addr_0}),
	.address_b({gnd,gnd,gnd,gnd,dc_tag_rd_port_addr_5,dc_tag_rd_port_addr_4,dc_tag_rd_port_addr_3,dc_tag_rd_port_addr_2,dc_tag_rd_port_addr_1,dc_tag_rd_port_addr_0}),
	.clock0(clk_clk));

endmodule

module embedded_system_altsyncram_3 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[9:0] address_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_v0o1 auto_generated(
	.q_b({q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.data_a({data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module embedded_system_altsyncram_v0o1 (
	q_b,
	wren_a,
	data_a,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[4:0] q_b;
input 	wren_a;
input 	[4:0] data_a;
input 	[5:0] address_a;
input 	[5:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "embedded_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_tag_module:embedded_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_v0o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 6;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 63;
defparam ram_block1a1.port_a_logical_ram_depth = 64;
defparam ram_block1a1.port_a_logical_ram_width = 5;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 6;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 63;
defparam ram_block1a1.port_b_logical_ram_depth = 64;
defparam ram_block1a1.port_b_logical_ram_width = 5;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "546805D71DAAEDDD";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "embedded_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_tag_module:embedded_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_v0o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 6;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 63;
defparam ram_block1a2.port_a_logical_ram_depth = 64;
defparam ram_block1a2.port_a_logical_ram_width = 5;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 6;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 63;
defparam ram_block1a2.port_b_logical_ram_depth = 64;
defparam ram_block1a2.port_b_logical_ram_width = 5;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "E2F31B031D14CD17";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "embedded_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_tag_module:embedded_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_v0o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 6;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 63;
defparam ram_block1a3.port_a_logical_ram_depth = 64;
defparam ram_block1a3.port_a_logical_ram_width = 5;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 6;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 63;
defparam ram_block1a3.port_b_logical_ram_depth = 64;
defparam ram_block1a3.port_b_logical_ram_width = 5;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "1F2ED13DF665EFF7";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "embedded_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_tag_module:embedded_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_v0o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 6;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 63;
defparam ram_block1a0.port_a_logical_ram_depth = 64;
defparam ram_block1a0.port_a_logical_ram_width = 5;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 6;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 63;
defparam ram_block1a0.port_b_logical_ram_depth = 64;
defparam ram_block1a0.port_b_logical_ram_width = 5;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "813B71E642DED444";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "embedded_system_nios2_qsys_0_dc_tag_ram.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_tag_module:embedded_system_nios2_qsys_0_dc_tag|altsyncram:the_altsyncram|altsyncram_v0o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 6;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 63;
defparam ram_block1a4.port_a_logical_ram_depth = 64;
defparam ram_block1a4.port_a_logical_ram_width = 5;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 6;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 63;
defparam ram_block1a4.port_b_logical_ram_depth = 64;
defparam ram_block1a4.port_b_logical_ram_width = 5;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "BC5E44A5DC51F506";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_dc_victim_module (
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_13,
	q_b_12,
	q_b_21,
	q_b_20,
	q_b_25,
	q_b_17,
	q_b_24,
	q_b_16,
	q_b_27,
	q_b_19,
	q_b_26,
	q_b_18,
	q_b_23,
	q_b_15,
	q_b_22,
	q_b_14,
	A_dc_xfer_wr_data_11,
	A_dc_xfer_wr_data_10,
	A_dc_xfer_wr_data_9,
	A_dc_xfer_wr_data_8,
	A_dc_xfer_wr_data_13,
	A_dc_xfer_wr_data_12,
	q_b_2,
	q_b_0,
	q_b_3,
	q_b_1,
	A_dc_xfer_wr_data_21,
	A_dc_xfer_wr_data_20,
	A_dc_xfer_wr_data_25,
	A_dc_xfer_wr_data_17,
	A_dc_xfer_wr_data_24,
	A_dc_xfer_wr_data_16,
	A_dc_xfer_wr_data_27,
	A_dc_xfer_wr_data_19,
	A_dc_xfer_wr_data_26,
	A_dc_xfer_wr_data_18,
	A_dc_xfer_wr_data_23,
	A_dc_xfer_wr_data_15,
	A_dc_xfer_wr_data_22,
	A_dc_xfer_wr_data_14,
	A_dc_xfer_wr_data_2,
	A_dc_xfer_wr_data_0,
	A_dc_xfer_wr_data_3,
	q_b_6,
	q_b_4,
	q_b_7,
	q_b_5,
	A_dc_xfer_wr_data_1,
	A_dc_xfer_wr_data_6,
	A_dc_xfer_wr_data_4,
	A_dc_xfer_wr_data_7,
	A_dc_xfer_wr_data_5,
	q_b_31,
	q_b_29,
	q_b_28,
	q_b_30,
	A_dc_xfer_wr_data_31,
	A_dc_xfer_wr_data_29,
	A_dc_xfer_wr_data_28,
	A_dc_xfer_wr_data_30,
	A_dc_xfer_wr_active,
	A_dc_wb_rd_en,
	A_dc_xfer_wr_offset_0,
	A_dc_xfer_wr_offset_1,
	A_dc_xfer_wr_offset_2,
	A_dc_wb_rd_addr_offset_0,
	A_dc_wb_rd_addr_offset_1,
	A_dc_wb_rd_addr_offset_2,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_13;
output 	q_b_12;
output 	q_b_21;
output 	q_b_20;
output 	q_b_25;
output 	q_b_17;
output 	q_b_24;
output 	q_b_16;
output 	q_b_27;
output 	q_b_19;
output 	q_b_26;
output 	q_b_18;
output 	q_b_23;
output 	q_b_15;
output 	q_b_22;
output 	q_b_14;
input 	A_dc_xfer_wr_data_11;
input 	A_dc_xfer_wr_data_10;
input 	A_dc_xfer_wr_data_9;
input 	A_dc_xfer_wr_data_8;
input 	A_dc_xfer_wr_data_13;
input 	A_dc_xfer_wr_data_12;
output 	q_b_2;
output 	q_b_0;
output 	q_b_3;
output 	q_b_1;
input 	A_dc_xfer_wr_data_21;
input 	A_dc_xfer_wr_data_20;
input 	A_dc_xfer_wr_data_25;
input 	A_dc_xfer_wr_data_17;
input 	A_dc_xfer_wr_data_24;
input 	A_dc_xfer_wr_data_16;
input 	A_dc_xfer_wr_data_27;
input 	A_dc_xfer_wr_data_19;
input 	A_dc_xfer_wr_data_26;
input 	A_dc_xfer_wr_data_18;
input 	A_dc_xfer_wr_data_23;
input 	A_dc_xfer_wr_data_15;
input 	A_dc_xfer_wr_data_22;
input 	A_dc_xfer_wr_data_14;
input 	A_dc_xfer_wr_data_2;
input 	A_dc_xfer_wr_data_0;
input 	A_dc_xfer_wr_data_3;
output 	q_b_6;
output 	q_b_4;
output 	q_b_7;
output 	q_b_5;
input 	A_dc_xfer_wr_data_1;
input 	A_dc_xfer_wr_data_6;
input 	A_dc_xfer_wr_data_4;
input 	A_dc_xfer_wr_data_7;
input 	A_dc_xfer_wr_data_5;
output 	q_b_31;
output 	q_b_29;
output 	q_b_28;
output 	q_b_30;
input 	A_dc_xfer_wr_data_31;
input 	A_dc_xfer_wr_data_29;
input 	A_dc_xfer_wr_data_28;
input 	A_dc_xfer_wr_data_30;
input 	A_dc_xfer_wr_active;
input 	A_dc_wb_rd_en;
input 	A_dc_xfer_wr_offset_0;
input 	A_dc_xfer_wr_offset_1;
input 	A_dc_xfer_wr_offset_2;
input 	A_dc_wb_rd_addr_offset_0;
input 	A_dc_wb_rd_addr_offset_1;
input 	A_dc_wb_rd_addr_offset_2;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_4 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({A_dc_xfer_wr_data_31,A_dc_xfer_wr_data_30,A_dc_xfer_wr_data_29,A_dc_xfer_wr_data_28,A_dc_xfer_wr_data_27,A_dc_xfer_wr_data_26,A_dc_xfer_wr_data_25,A_dc_xfer_wr_data_24,A_dc_xfer_wr_data_23,A_dc_xfer_wr_data_22,A_dc_xfer_wr_data_21,A_dc_xfer_wr_data_20,
A_dc_xfer_wr_data_19,A_dc_xfer_wr_data_18,A_dc_xfer_wr_data_17,A_dc_xfer_wr_data_16,A_dc_xfer_wr_data_15,A_dc_xfer_wr_data_14,A_dc_xfer_wr_data_13,A_dc_xfer_wr_data_12,A_dc_xfer_wr_data_11,A_dc_xfer_wr_data_10,A_dc_xfer_wr_data_9,A_dc_xfer_wr_data_8,
A_dc_xfer_wr_data_7,A_dc_xfer_wr_data_6,A_dc_xfer_wr_data_5,A_dc_xfer_wr_data_4,A_dc_xfer_wr_data_3,A_dc_xfer_wr_data_2,A_dc_xfer_wr_data_1,A_dc_xfer_wr_data_0}),
	.wren_a(A_dc_xfer_wr_active),
	.rden_b(A_dc_wb_rd_en),
	.address_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_dc_xfer_wr_offset_2,A_dc_xfer_wr_offset_1,A_dc_xfer_wr_offset_0}),
	.address_b({gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_dc_wb_rd_addr_offset_2,A_dc_wb_rd_addr_offset_1,A_dc_wb_rd_addr_offset_0}),
	.clock0(clk_clk));

endmodule

module embedded_system_altsyncram_4 (
	q_b,
	data_a,
	wren_a,
	rden_b,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	wren_a;
input 	rden_b;
input 	[9:0] address_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_baj1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.wren_a(wren_a),
	.rden_b(rden_b),
	.address_a({address_a[2],address_a[1],address_a[0]}),
	.address_b({address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module embedded_system_altsyncram_baj1 (
	q_b,
	data_a,
	wren_a,
	rden_b,
	address_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	wren_a;
input 	rden_b;
input 	[2:0] address_a;
input 	[2:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 3;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 7;
defparam ram_block1a11.port_a_logical_ram_depth = 8;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 3;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 7;
defparam ram_block1a11.port_b_logical_ram_depth = 8;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 3;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 7;
defparam ram_block1a10.port_a_logical_ram_depth = 8;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 3;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 7;
defparam ram_block1a10.port_b_logical_ram_depth = 8;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 3;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 7;
defparam ram_block1a9.port_a_logical_ram_depth = 8;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 3;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 7;
defparam ram_block1a9.port_b_logical_ram_depth = 8;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 3;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 7;
defparam ram_block1a8.port_a_logical_ram_depth = 8;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 3;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 7;
defparam ram_block1a13.port_a_logical_ram_depth = 8;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 3;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 7;
defparam ram_block1a13.port_b_logical_ram_depth = 8;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 3;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 7;
defparam ram_block1a12.port_a_logical_ram_depth = 8;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 3;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 7;
defparam ram_block1a12.port_b_logical_ram_depth = 8;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 3;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 7;
defparam ram_block1a21.port_a_logical_ram_depth = 8;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 3;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 7;
defparam ram_block1a21.port_b_logical_ram_depth = 8;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 3;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 7;
defparam ram_block1a20.port_a_logical_ram_depth = 8;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 3;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 7;
defparam ram_block1a20.port_b_logical_ram_depth = 8;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 3;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 7;
defparam ram_block1a25.port_a_logical_ram_depth = 8;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 3;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 7;
defparam ram_block1a25.port_b_logical_ram_depth = 8;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 3;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 7;
defparam ram_block1a17.port_a_logical_ram_depth = 8;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 3;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 7;
defparam ram_block1a17.port_b_logical_ram_depth = 8;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 3;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 7;
defparam ram_block1a24.port_a_logical_ram_depth = 8;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 3;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 7;
defparam ram_block1a24.port_b_logical_ram_depth = 8;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 3;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 7;
defparam ram_block1a16.port_a_logical_ram_depth = 8;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 3;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 7;
defparam ram_block1a16.port_b_logical_ram_depth = 8;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 3;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 7;
defparam ram_block1a27.port_a_logical_ram_depth = 8;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 3;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 7;
defparam ram_block1a27.port_b_logical_ram_depth = 8;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 3;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 7;
defparam ram_block1a19.port_a_logical_ram_depth = 8;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 3;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 7;
defparam ram_block1a19.port_b_logical_ram_depth = 8;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 3;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 7;
defparam ram_block1a26.port_a_logical_ram_depth = 8;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 3;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 7;
defparam ram_block1a26.port_b_logical_ram_depth = 8;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 3;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 7;
defparam ram_block1a18.port_a_logical_ram_depth = 8;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 3;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 7;
defparam ram_block1a18.port_b_logical_ram_depth = 8;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 3;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 7;
defparam ram_block1a23.port_a_logical_ram_depth = 8;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 3;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 7;
defparam ram_block1a23.port_b_logical_ram_depth = 8;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 3;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 7;
defparam ram_block1a15.port_a_logical_ram_depth = 8;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 3;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 7;
defparam ram_block1a15.port_b_logical_ram_depth = 8;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 3;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 7;
defparam ram_block1a22.port_a_logical_ram_depth = 8;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 3;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 7;
defparam ram_block1a22.port_b_logical_ram_depth = 8;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 3;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 7;
defparam ram_block1a14.port_a_logical_ram_depth = 8;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 3;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 7;
defparam ram_block1a14.port_b_logical_ram_depth = 8;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 3;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 7;
defparam ram_block1a2.port_a_logical_ram_depth = 8;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 3;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 7;
defparam ram_block1a2.port_b_logical_ram_depth = 8;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 3;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 7;
defparam ram_block1a0.port_a_logical_ram_depth = 8;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 3;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 7;
defparam ram_block1a0.port_b_logical_ram_depth = 8;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 3;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 7;
defparam ram_block1a3.port_a_logical_ram_depth = 8;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 3;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 7;
defparam ram_block1a3.port_b_logical_ram_depth = 8;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 3;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 7;
defparam ram_block1a1.port_a_logical_ram_depth = 8;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 3;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 7;
defparam ram_block1a1.port_b_logical_ram_depth = 8;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 3;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 7;
defparam ram_block1a6.port_a_logical_ram_depth = 8;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 3;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 7;
defparam ram_block1a4.port_a_logical_ram_depth = 8;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 3;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 7;
defparam ram_block1a7.port_a_logical_ram_depth = 8;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 3;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 7;
defparam ram_block1a5.port_a_logical_ram_depth = 8;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 3;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 7;
defparam ram_block1a31.port_a_logical_ram_depth = 8;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 3;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 7;
defparam ram_block1a31.port_b_logical_ram_depth = 8;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 3;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 7;
defparam ram_block1a29.port_a_logical_ram_depth = 8;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 3;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 7;
defparam ram_block1a29.port_b_logical_ram_depth = 8;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 3;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 7;
defparam ram_block1a28.port_a_logical_ram_depth = 8;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 3;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 7;
defparam ram_block1a28.port_b_logical_ram_depth = 8;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_dc_victim_module:embedded_system_nios2_qsys_0_dc_victim|altsyncram:the_altsyncram|altsyncram_baj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 3;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 7;
defparam ram_block1a30.port_a_logical_ram_depth = 8;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 3;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 7;
defparam ram_block1a30.port_b_logical_ram_depth = 8;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_ic_data_module (
	q_b_5,
	q_b_3,
	q_b_1,
	q_b_4,
	q_b_2,
	q_b_28,
	q_b_31,
	q_b_27,
	q_b_29,
	q_b_30,
	q_b_0,
	q_b_23,
	q_b_26,
	q_b_22,
	q_b_24,
	q_b_25,
	q_b_16,
	q_b_15,
	q_b_13,
	q_b_14,
	q_b_12,
	q_b_11,
	q_b_8,
	q_b_19,
	q_b_18,
	q_b_17,
	q_b_10,
	q_b_9,
	q_b_21,
	q_b_20,
	q_b_7,
	q_b_6,
	ic_fill_line_6,
	ic_fill_line_5,
	ic_fill_line_1,
	ic_fill_line_0,
	ic_fill_line_4,
	ic_fill_line_3,
	ic_fill_line_2,
	F_stall,
	ic_fill_dp_offset_0,
	ic_fill_dp_offset_1,
	ic_fill_dp_offset_2,
	i_readdatavalid_d1,
	i_readdata_d1_5,
	F_ic_data_rd_addr_nxt_0,
	F_ic_data_rd_addr_nxt_1,
	F_ic_data_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_0,
	F_ic_tag_rd_addr_nxt_1,
	F_ic_tag_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_3,
	F_ic_tag_rd_addr_nxt_4,
	F_ic_tag_rd_addr_nxt_5,
	F_ic_tag_rd_addr_nxt_6,
	i_readdata_d1_3,
	i_readdata_d1_1,
	i_readdata_d1_4,
	i_readdata_d1_2,
	i_readdata_d1_28,
	i_readdata_d1_31,
	i_readdata_d1_27,
	i_readdata_d1_29,
	i_readdata_d1_30,
	i_readdata_d1_0,
	i_readdata_d1_23,
	i_readdata_d1_26,
	i_readdata_d1_22,
	i_readdata_d1_24,
	i_readdata_d1_25,
	i_readdata_d1_16,
	i_readdata_d1_15,
	i_readdata_d1_13,
	i_readdata_d1_14,
	i_readdata_d1_12,
	i_readdata_d1_11,
	i_readdata_d1_8,
	i_readdata_d1_19,
	i_readdata_d1_18,
	i_readdata_d1_17,
	i_readdata_d1_10,
	i_readdata_d1_9,
	i_readdata_d1_21,
	i_readdata_d1_20,
	i_readdata_d1_7,
	i_readdata_d1_6,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_5;
output 	q_b_3;
output 	q_b_1;
output 	q_b_4;
output 	q_b_2;
output 	q_b_28;
output 	q_b_31;
output 	q_b_27;
output 	q_b_29;
output 	q_b_30;
output 	q_b_0;
output 	q_b_23;
output 	q_b_26;
output 	q_b_22;
output 	q_b_24;
output 	q_b_25;
output 	q_b_16;
output 	q_b_15;
output 	q_b_13;
output 	q_b_14;
output 	q_b_12;
output 	q_b_11;
output 	q_b_8;
output 	q_b_19;
output 	q_b_18;
output 	q_b_17;
output 	q_b_10;
output 	q_b_9;
output 	q_b_21;
output 	q_b_20;
output 	q_b_7;
output 	q_b_6;
input 	ic_fill_line_6;
input 	ic_fill_line_5;
input 	ic_fill_line_1;
input 	ic_fill_line_0;
input 	ic_fill_line_4;
input 	ic_fill_line_3;
input 	ic_fill_line_2;
input 	F_stall;
input 	ic_fill_dp_offset_0;
input 	ic_fill_dp_offset_1;
input 	ic_fill_dp_offset_2;
input 	i_readdatavalid_d1;
input 	i_readdata_d1_5;
input 	F_ic_data_rd_addr_nxt_0;
input 	F_ic_data_rd_addr_nxt_1;
input 	F_ic_data_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_0;
input 	F_ic_tag_rd_addr_nxt_1;
input 	F_ic_tag_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_3;
input 	F_ic_tag_rd_addr_nxt_4;
input 	F_ic_tag_rd_addr_nxt_5;
input 	F_ic_tag_rd_addr_nxt_6;
input 	i_readdata_d1_3;
input 	i_readdata_d1_1;
input 	i_readdata_d1_4;
input 	i_readdata_d1_2;
input 	i_readdata_d1_28;
input 	i_readdata_d1_31;
input 	i_readdata_d1_27;
input 	i_readdata_d1_29;
input 	i_readdata_d1_30;
input 	i_readdata_d1_0;
input 	i_readdata_d1_23;
input 	i_readdata_d1_26;
input 	i_readdata_d1_22;
input 	i_readdata_d1_24;
input 	i_readdata_d1_25;
input 	i_readdata_d1_16;
input 	i_readdata_d1_15;
input 	i_readdata_d1_13;
input 	i_readdata_d1_14;
input 	i_readdata_d1_12;
input 	i_readdata_d1_11;
input 	i_readdata_d1_8;
input 	i_readdata_d1_19;
input 	i_readdata_d1_18;
input 	i_readdata_d1_17;
input 	i_readdata_d1_10;
input 	i_readdata_d1_9;
input 	i_readdata_d1_21;
input 	i_readdata_d1_20;
input 	i_readdata_d1_7;
input 	i_readdata_d1_6;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_5 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({ic_fill_line_6,ic_fill_line_5,ic_fill_line_4,ic_fill_line_3,ic_fill_line_2,ic_fill_line_1,ic_fill_line_0,ic_fill_dp_offset_2,ic_fill_dp_offset_1,ic_fill_dp_offset_0}),
	.rden_b(F_stall),
	.wren_a(i_readdatavalid_d1),
	.data_a({i_readdata_d1_31,i_readdata_d1_30,i_readdata_d1_29,i_readdata_d1_28,i_readdata_d1_27,i_readdata_d1_26,i_readdata_d1_25,i_readdata_d1_24,i_readdata_d1_23,i_readdata_d1_22,i_readdata_d1_21,i_readdata_d1_20,i_readdata_d1_19,i_readdata_d1_18,i_readdata_d1_17,i_readdata_d1_16,
i_readdata_d1_15,i_readdata_d1_14,i_readdata_d1_13,i_readdata_d1_12,i_readdata_d1_11,i_readdata_d1_10,i_readdata_d1_9,i_readdata_d1_8,i_readdata_d1_7,i_readdata_d1_6,i_readdata_d1_5,i_readdata_d1_4,i_readdata_d1_3,i_readdata_d1_2,i_readdata_d1_1,i_readdata_d1_0}),
	.address_b({F_ic_tag_rd_addr_nxt_6,F_ic_tag_rd_addr_nxt_5,F_ic_tag_rd_addr_nxt_4,F_ic_tag_rd_addr_nxt_3,F_ic_tag_rd_addr_nxt_2,F_ic_tag_rd_addr_nxt_1,F_ic_tag_rd_addr_nxt_0,F_ic_data_rd_addr_nxt_2,F_ic_data_rd_addr_nxt_1,F_ic_data_rd_addr_nxt_0}),
	.clock0(clk_clk));

endmodule

module embedded_system_altsyncram_5 (
	q_b,
	address_a,
	rden_b,
	wren_a,
	data_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[9:0] address_a;
input 	rden_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_spj1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.rden_b(rden_b),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_b({address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module embedded_system_altsyncram_spj1 (
	q_b,
	address_a,
	rden_b,
	wren_a,
	data_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[9:0] address_a;
input 	rden_b;
input 	wren_a;
input 	[31:0] data_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk1_core_clock_enable = "ena1";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 10;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 1023;
defparam ram_block1a5.port_a_logical_ram_depth = 1024;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock1";
defparam ram_block1a5.port_b_address_width = 10;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 1023;
defparam ram_block1a5.port_b_logical_ram_depth = 1024;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock1";
defparam ram_block1a5.ram_block_type = "auto";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk1_core_clock_enable = "ena1";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 10;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 1023;
defparam ram_block1a3.port_a_logical_ram_depth = 1024;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock1";
defparam ram_block1a3.port_b_address_width = 10;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 1023;
defparam ram_block1a3.port_b_logical_ram_depth = 1024;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock1";
defparam ram_block1a3.ram_block_type = "auto";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk1_core_clock_enable = "ena1";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 10;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 1023;
defparam ram_block1a1.port_a_logical_ram_depth = 1024;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock1";
defparam ram_block1a1.port_b_address_width = 10;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 1023;
defparam ram_block1a1.port_b_logical_ram_depth = 1024;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock1";
defparam ram_block1a1.ram_block_type = "auto";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk1_core_clock_enable = "ena1";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 10;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 1023;
defparam ram_block1a4.port_a_logical_ram_depth = 1024;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock1";
defparam ram_block1a4.port_b_address_width = 10;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 1023;
defparam ram_block1a4.port_b_logical_ram_depth = 1024;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock1";
defparam ram_block1a4.ram_block_type = "auto";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk1_core_clock_enable = "ena1";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 10;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 1023;
defparam ram_block1a2.port_a_logical_ram_depth = 1024;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock1";
defparam ram_block1a2.port_b_address_width = 10;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 1023;
defparam ram_block1a2.port_b_logical_ram_depth = 1024;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock1";
defparam ram_block1a2.ram_block_type = "auto";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk1_core_clock_enable = "ena1";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 10;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 1023;
defparam ram_block1a28.port_a_logical_ram_depth = 1024;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock1";
defparam ram_block1a28.port_b_address_width = 10;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 1023;
defparam ram_block1a28.port_b_logical_ram_depth = 1024;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock1";
defparam ram_block1a28.ram_block_type = "auto";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk1_core_clock_enable = "ena1";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 10;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 1023;
defparam ram_block1a31.port_a_logical_ram_depth = 1024;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock1";
defparam ram_block1a31.port_b_address_width = 10;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 1023;
defparam ram_block1a31.port_b_logical_ram_depth = 1024;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock1";
defparam ram_block1a31.ram_block_type = "auto";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk1_core_clock_enable = "ena1";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 10;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 1023;
defparam ram_block1a27.port_a_logical_ram_depth = 1024;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock1";
defparam ram_block1a27.port_b_address_width = 10;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 1023;
defparam ram_block1a27.port_b_logical_ram_depth = 1024;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock1";
defparam ram_block1a27.ram_block_type = "auto";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk1_core_clock_enable = "ena1";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 10;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 1023;
defparam ram_block1a29.port_a_logical_ram_depth = 1024;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock1";
defparam ram_block1a29.port_b_address_width = 10;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 1023;
defparam ram_block1a29.port_b_logical_ram_depth = 1024;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock1";
defparam ram_block1a29.ram_block_type = "auto";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk1_core_clock_enable = "ena1";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 10;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 1023;
defparam ram_block1a30.port_a_logical_ram_depth = 1024;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock1";
defparam ram_block1a30.port_b_address_width = 10;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 1023;
defparam ram_block1a30.port_b_logical_ram_depth = 1024;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock1";
defparam ram_block1a30.ram_block_type = "auto";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk1_core_clock_enable = "ena1";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 10;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 1023;
defparam ram_block1a0.port_a_logical_ram_depth = 1024;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock1";
defparam ram_block1a0.port_b_address_width = 10;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 1023;
defparam ram_block1a0.port_b_logical_ram_depth = 1024;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock1";
defparam ram_block1a0.ram_block_type = "auto";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk1_core_clock_enable = "ena1";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 10;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 1023;
defparam ram_block1a23.port_a_logical_ram_depth = 1024;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock1";
defparam ram_block1a23.port_b_address_width = 10;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 1023;
defparam ram_block1a23.port_b_logical_ram_depth = 1024;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock1";
defparam ram_block1a23.ram_block_type = "auto";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk1_core_clock_enable = "ena1";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 10;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 1023;
defparam ram_block1a26.port_a_logical_ram_depth = 1024;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock1";
defparam ram_block1a26.port_b_address_width = 10;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 1023;
defparam ram_block1a26.port_b_logical_ram_depth = 1024;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock1";
defparam ram_block1a26.ram_block_type = "auto";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk1_core_clock_enable = "ena1";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 10;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 1023;
defparam ram_block1a22.port_a_logical_ram_depth = 1024;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock1";
defparam ram_block1a22.port_b_address_width = 10;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 1023;
defparam ram_block1a22.port_b_logical_ram_depth = 1024;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock1";
defparam ram_block1a22.ram_block_type = "auto";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk1_core_clock_enable = "ena1";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 10;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 1023;
defparam ram_block1a24.port_a_logical_ram_depth = 1024;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock1";
defparam ram_block1a24.port_b_address_width = 10;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 1023;
defparam ram_block1a24.port_b_logical_ram_depth = 1024;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock1";
defparam ram_block1a24.ram_block_type = "auto";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk1_core_clock_enable = "ena1";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 10;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 1023;
defparam ram_block1a25.port_a_logical_ram_depth = 1024;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock1";
defparam ram_block1a25.port_b_address_width = 10;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 1023;
defparam ram_block1a25.port_b_logical_ram_depth = 1024;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock1";
defparam ram_block1a25.ram_block_type = "auto";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk1_core_clock_enable = "ena1";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 10;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 1023;
defparam ram_block1a16.port_a_logical_ram_depth = 1024;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock1";
defparam ram_block1a16.port_b_address_width = 10;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 1023;
defparam ram_block1a16.port_b_logical_ram_depth = 1024;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock1";
defparam ram_block1a16.ram_block_type = "auto";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk1_core_clock_enable = "ena1";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 10;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 1023;
defparam ram_block1a15.port_a_logical_ram_depth = 1024;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock1";
defparam ram_block1a15.port_b_address_width = 10;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 1023;
defparam ram_block1a15.port_b_logical_ram_depth = 1024;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock1";
defparam ram_block1a15.ram_block_type = "auto";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk1_core_clock_enable = "ena1";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 10;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 1023;
defparam ram_block1a13.port_a_logical_ram_depth = 1024;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock1";
defparam ram_block1a13.port_b_address_width = 10;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 1023;
defparam ram_block1a13.port_b_logical_ram_depth = 1024;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock1";
defparam ram_block1a13.ram_block_type = "auto";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk1_core_clock_enable = "ena1";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 10;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 1023;
defparam ram_block1a14.port_a_logical_ram_depth = 1024;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock1";
defparam ram_block1a14.port_b_address_width = 10;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 1023;
defparam ram_block1a14.port_b_logical_ram_depth = 1024;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock1";
defparam ram_block1a14.ram_block_type = "auto";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk1_core_clock_enable = "ena1";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 10;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 1023;
defparam ram_block1a12.port_a_logical_ram_depth = 1024;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock1";
defparam ram_block1a12.port_b_address_width = 10;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 1023;
defparam ram_block1a12.port_b_logical_ram_depth = 1024;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock1";
defparam ram_block1a12.ram_block_type = "auto";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk1_core_clock_enable = "ena1";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 10;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 1023;
defparam ram_block1a11.port_a_logical_ram_depth = 1024;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock1";
defparam ram_block1a11.port_b_address_width = 10;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 1023;
defparam ram_block1a11.port_b_logical_ram_depth = 1024;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock1";
defparam ram_block1a11.ram_block_type = "auto";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk1_core_clock_enable = "ena1";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 10;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 1023;
defparam ram_block1a8.port_a_logical_ram_depth = 1024;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock1";
defparam ram_block1a8.port_b_address_width = 10;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 1023;
defparam ram_block1a8.port_b_logical_ram_depth = 1024;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock1";
defparam ram_block1a8.ram_block_type = "auto";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk1_core_clock_enable = "ena1";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 10;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 1023;
defparam ram_block1a19.port_a_logical_ram_depth = 1024;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock1";
defparam ram_block1a19.port_b_address_width = 10;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 1023;
defparam ram_block1a19.port_b_logical_ram_depth = 1024;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock1";
defparam ram_block1a19.ram_block_type = "auto";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk1_core_clock_enable = "ena1";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 10;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 1023;
defparam ram_block1a18.port_a_logical_ram_depth = 1024;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock1";
defparam ram_block1a18.port_b_address_width = 10;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 1023;
defparam ram_block1a18.port_b_logical_ram_depth = 1024;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock1";
defparam ram_block1a18.ram_block_type = "auto";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk1_core_clock_enable = "ena1";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 10;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 1023;
defparam ram_block1a17.port_a_logical_ram_depth = 1024;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock1";
defparam ram_block1a17.port_b_address_width = 10;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 1023;
defparam ram_block1a17.port_b_logical_ram_depth = 1024;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock1";
defparam ram_block1a17.ram_block_type = "auto";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk1_core_clock_enable = "ena1";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 10;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 1023;
defparam ram_block1a10.port_a_logical_ram_depth = 1024;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock1";
defparam ram_block1a10.port_b_address_width = 10;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 1023;
defparam ram_block1a10.port_b_logical_ram_depth = 1024;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock1";
defparam ram_block1a10.ram_block_type = "auto";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk1_core_clock_enable = "ena1";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 10;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 1023;
defparam ram_block1a9.port_a_logical_ram_depth = 1024;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock1";
defparam ram_block1a9.port_b_address_width = 10;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 1023;
defparam ram_block1a9.port_b_logical_ram_depth = 1024;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock1";
defparam ram_block1a9.ram_block_type = "auto";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk1_core_clock_enable = "ena1";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 10;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 1023;
defparam ram_block1a21.port_a_logical_ram_depth = 1024;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock1";
defparam ram_block1a21.port_b_address_width = 10;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 1023;
defparam ram_block1a21.port_b_logical_ram_depth = 1024;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock1";
defparam ram_block1a21.ram_block_type = "auto";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk1_core_clock_enable = "ena1";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 10;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 1023;
defparam ram_block1a20.port_a_logical_ram_depth = 1024;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock1";
defparam ram_block1a20.port_b_address_width = 10;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 1023;
defparam ram_block1a20.port_b_logical_ram_depth = 1024;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock1";
defparam ram_block1a20.ram_block_type = "auto";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk1_core_clock_enable = "ena1";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 10;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 1023;
defparam ram_block1a7.port_a_logical_ram_depth = 1024;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock1";
defparam ram_block1a7.port_b_address_width = 10;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 1023;
defparam ram_block1a7.port_b_logical_ram_depth = 1024;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock1";
defparam ram_block1a7.ram_block_type = "auto";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock0),
	.ena0(wren_a),
	.ena1(!rden_b),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk1_core_clock_enable = "ena1";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_data_module:embedded_system_nios2_qsys_0_ic_data|altsyncram:the_altsyncram|altsyncram_spj1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 10;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 1023;
defparam ram_block1a6.port_a_logical_ram_depth = 1024;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock1";
defparam ram_block1a6.port_b_address_width = 10;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 1023;
defparam ram_block1a6.port_b_logical_ram_depth = 1024;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock1";
defparam ram_block1a6.ram_block_type = "auto";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_ic_tag_module (
	q_b_0,
	q_b_1,
	q_b_7,
	q_b_9,
	q_b_6,
	q_b_8,
	ic_fill_valid_bits_5,
	ic_fill_valid_bits_7,
	ic_fill_valid_bits_4,
	q_b_3,
	q_b_5,
	q_b_2,
	q_b_4,
	ic_fill_valid_bits_6,
	ic_fill_valid_bits_1,
	ic_fill_valid_bits_3,
	ic_fill_valid_bits_0,
	ic_fill_valid_bits_2,
	ic_fill_tag_1,
	ic_fill_tag_0,
	F_stall,
	F_ic_tag_rd_addr_nxt_0,
	F_ic_tag_rd_addr_nxt_1,
	F_ic_tag_rd_addr_nxt_2,
	F_ic_tag_rd_addr_nxt_3,
	F_ic_tag_rd_addr_nxt_4,
	F_ic_tag_rd_addr_nxt_5,
	F_ic_tag_rd_addr_nxt_6,
	ic_tag_wren,
	ic_tag_wraddress_0,
	ic_tag_wraddress_1,
	ic_tag_wraddress_2,
	ic_tag_wraddress_3,
	ic_tag_wraddress_4,
	ic_tag_wraddress_5,
	ic_tag_wraddress_6,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_0;
output 	q_b_1;
output 	q_b_7;
output 	q_b_9;
output 	q_b_6;
output 	q_b_8;
input 	ic_fill_valid_bits_5;
input 	ic_fill_valid_bits_7;
input 	ic_fill_valid_bits_4;
output 	q_b_3;
output 	q_b_5;
output 	q_b_2;
output 	q_b_4;
input 	ic_fill_valid_bits_6;
input 	ic_fill_valid_bits_1;
input 	ic_fill_valid_bits_3;
input 	ic_fill_valid_bits_0;
input 	ic_fill_valid_bits_2;
input 	ic_fill_tag_1;
input 	ic_fill_tag_0;
input 	F_stall;
input 	F_ic_tag_rd_addr_nxt_0;
input 	F_ic_tag_rd_addr_nxt_1;
input 	F_ic_tag_rd_addr_nxt_2;
input 	F_ic_tag_rd_addr_nxt_3;
input 	F_ic_tag_rd_addr_nxt_4;
input 	F_ic_tag_rd_addr_nxt_5;
input 	F_ic_tag_rd_addr_nxt_6;
input 	ic_tag_wren;
input 	ic_tag_wraddress_0;
input 	ic_tag_wraddress_1;
input 	ic_tag_wraddress_2;
input 	ic_tag_wraddress_3;
input 	ic_tag_wraddress_4;
input 	ic_tag_wraddress_5;
input 	ic_tag_wraddress_6;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_6 the_altsyncram(
	.q_b({q_b_unconnected_wire_31,q_b_unconnected_wire_30,q_b_unconnected_wire_29,q_b_unconnected_wire_28,q_b_unconnected_wire_27,q_b_unconnected_wire_26,q_b_unconnected_wire_25,q_b_unconnected_wire_24,q_b_unconnected_wire_23,q_b_unconnected_wire_22,q_b_unconnected_wire_21,
q_b_unconnected_wire_20,q_b_unconnected_wire_19,q_b_unconnected_wire_18,q_b_unconnected_wire_17,q_b_unconnected_wire_16,q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,
q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,ic_fill_valid_bits_7,ic_fill_valid_bits_6,ic_fill_valid_bits_5,ic_fill_valid_bits_4,ic_fill_valid_bits_3,ic_fill_valid_bits_2,ic_fill_valid_bits_1,ic_fill_valid_bits_0,ic_fill_tag_1,ic_fill_tag_0}),
	.rden_b(F_stall),
	.address_b({gnd,gnd,gnd,F_ic_tag_rd_addr_nxt_6,F_ic_tag_rd_addr_nxt_5,F_ic_tag_rd_addr_nxt_4,F_ic_tag_rd_addr_nxt_3,F_ic_tag_rd_addr_nxt_2,F_ic_tag_rd_addr_nxt_1,F_ic_tag_rd_addr_nxt_0}),
	.wren_a(ic_tag_wren),
	.address_a({gnd,gnd,gnd,ic_tag_wraddress_6,ic_tag_wraddress_5,ic_tag_wraddress_4,ic_tag_wraddress_3,ic_tag_wraddress_2,ic_tag_wraddress_1,ic_tag_wraddress_0}),
	.clock0(clk_clk));

endmodule

module embedded_system_altsyncram_6 (
	q_b,
	data_a,
	rden_b,
	address_b,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	rden_b;
input 	[9:0] address_b;
input 	wren_a;
input 	[9:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_aro1 auto_generated(
	.q_b({q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.rden_b(rden_b),
	.address_b({address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.wren_a(wren_a),
	.address_a({address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.clock0(clock0));

endmodule

module embedded_system_altsyncram_aro1 (
	q_b,
	data_a,
	rden_b,
	address_b,
	wren_a,
	address_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[9:0] q_b;
input 	[9:0] data_a;
input 	rden_b;
input 	[6:0] address_b;
input 	wren_a;
input 	[6:0] address_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "embedded_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_tag_module:embedded_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_aro1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 7;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 127;
defparam ram_block1a0.port_a_logical_ram_depth = 128;
defparam ram_block1a0.port_a_logical_ram_width = 10;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 7;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 127;
defparam ram_block1a0.port_b_logical_ram_depth = 128;
defparam ram_block1a0.port_b_logical_ram_width = 10;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "94A9F5690E3630A78C8585FC4B85E2D1";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "embedded_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_tag_module:embedded_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_aro1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 7;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 127;
defparam ram_block1a1.port_a_logical_ram_depth = 128;
defparam ram_block1a1.port_a_logical_ram_width = 10;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 7;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 127;
defparam ram_block1a1.port_b_logical_ram_depth = 128;
defparam ram_block1a1.port_b_logical_ram_width = 10;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "EDA981B22281FC5F11F642ED9054AB2E";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "embedded_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a7.init_file_layout = "port_b";
defparam ram_block1a7.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_tag_module:embedded_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_aro1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 7;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 127;
defparam ram_block1a7.port_a_logical_ram_depth = 128;
defparam ram_block1a7.port_a_logical_ram_width = 10;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 7;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 127;
defparam ram_block1a7.port_b_logical_ram_depth = 128;
defparam ram_block1a7.port_b_logical_ram_width = 10;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "655AED0BDD5E17898E90410A92DC1ACD";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "embedded_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a9.init_file_layout = "port_b";
defparam ram_block1a9.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_tag_module:embedded_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_aro1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 7;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 127;
defparam ram_block1a9.port_a_logical_ram_depth = 128;
defparam ram_block1a9.port_a_logical_ram_width = 10;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 7;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 127;
defparam ram_block1a9.port_b_logical_ram_depth = 128;
defparam ram_block1a9.port_b_logical_ram_width = 10;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "8801DDD5C912235A1E8A083C13FBB55F";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "embedded_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a6.init_file_layout = "port_b";
defparam ram_block1a6.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_tag_module:embedded_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_aro1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 7;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 127;
defparam ram_block1a6.port_a_logical_ram_depth = 128;
defparam ram_block1a6.port_a_logical_ram_width = 10;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 7;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 127;
defparam ram_block1a6.port_b_logical_ram_depth = 128;
defparam ram_block1a6.port_b_logical_ram_width = 10;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "658EBF19163FDCF68B8CE62A381885D2";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "embedded_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a8.init_file_layout = "port_b";
defparam ram_block1a8.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_tag_module:embedded_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_aro1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 7;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 127;
defparam ram_block1a8.port_a_logical_ram_depth = 128;
defparam ram_block1a8.port_a_logical_ram_width = 10;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 7;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 127;
defparam ram_block1a8.port_b_logical_ram_depth = 128;
defparam ram_block1a8.port_b_logical_ram_width = 10;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "5E7F197F35D17B123B1B82F59E89CCF4";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "embedded_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_tag_module:embedded_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_aro1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 7;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 127;
defparam ram_block1a3.port_a_logical_ram_depth = 128;
defparam ram_block1a3.port_a_logical_ram_width = 10;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 7;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 127;
defparam ram_block1a3.port_b_logical_ram_depth = 128;
defparam ram_block1a3.port_b_logical_ram_width = 10;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "0943CB764E2420468D3B27532E65E41F";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "embedded_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a5.init_file_layout = "port_b";
defparam ram_block1a5.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_tag_module:embedded_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_aro1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 7;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 127;
defparam ram_block1a5.port_a_logical_ram_depth = 128;
defparam ram_block1a5.port_a_logical_ram_width = 10;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 7;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 127;
defparam ram_block1a5.port_b_logical_ram_depth = 128;
defparam ram_block1a5.port_b_logical_ram_width = 10;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "0E43F1BDDE880511A2F0C3183652592A";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "embedded_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_tag_module:embedded_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_aro1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 7;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 127;
defparam ram_block1a2.port_a_logical_ram_depth = 128;
defparam ram_block1a2.port_a_logical_ram_width = 10;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 7;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 127;
defparam ram_block1a2.port_b_logical_ram_depth = 128;
defparam ram_block1a2.port_b_logical_ram_width = 10;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "09331835E02E36B16F157A2C9AA14D00";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(!rden_b),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "embedded_system_nios2_qsys_0_ic_tag_ram.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_ic_tag_module:embedded_system_nios2_qsys_0_ic_tag|altsyncram:the_altsyncram|altsyncram_aro1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 7;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 127;
defparam ram_block1a4.port_a_logical_ram_depth = 128;
defparam ram_block1a4.port_a_logical_ram_width = 10;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 7;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 127;
defparam ram_block1a4.port_b_logical_ram_depth = 128;
defparam ram_block1a4.port_b_logical_ram_width = 10;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "5C0AC6C6BC7F5E1D56C5C85B156BC2F6";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_mult_cell (
	Add0,
	Add01,
	Add02,
	Add03,
	Add04,
	Add05,
	Add06,
	Add07,
	Add08,
	Add09,
	Add010,
	Add011,
	Add012,
	Add013,
	Add014,
	Add015,
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_0,
	A_mul_src1_1,
	A_mul_src1_2,
	A_mul_src1_3,
	A_mul_src1_4,
	A_mul_src1_5,
	A_mul_src1_6,
	A_mul_src1_7,
	A_mul_src1_8,
	A_mul_src1_9,
	A_mul_src1_10,
	A_mul_src1_11,
	A_mul_src1_12,
	A_mul_src1_13,
	A_mul_src1_14,
	A_mul_src1_15,
	A_mul_src1_16,
	A_mul_src1_17,
	A_mul_src1_18,
	A_mul_src1_19,
	A_mul_src1_20,
	A_mul_src1_21,
	A_mul_src1_22,
	A_mul_src1_23,
	A_mul_src1_24,
	A_mul_src1_25,
	A_mul_src1_26,
	A_mul_src1_27,
	A_mul_src1_28,
	A_mul_src1_29,
	A_mul_src1_30,
	A_mul_src1_31,
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	data_out_wire_2,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_0,
	data_out_wire_15,
	data_out_wire_14,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	Add0;
output 	Add01;
output 	Add02;
output 	Add03;
output 	Add04;
output 	Add05;
output 	Add06;
output 	Add07;
output 	Add08;
output 	Add09;
output 	Add010;
output 	Add011;
output 	Add012;
output 	Add013;
output 	Add014;
output 	Add015;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_0;
input 	A_mul_src1_1;
input 	A_mul_src1_2;
input 	A_mul_src1_3;
input 	A_mul_src1_4;
input 	A_mul_src1_5;
input 	A_mul_src1_6;
input 	A_mul_src1_7;
input 	A_mul_src1_8;
input 	A_mul_src1_9;
input 	A_mul_src1_10;
input 	A_mul_src1_11;
input 	A_mul_src1_12;
input 	A_mul_src1_13;
input 	A_mul_src1_14;
input 	A_mul_src1_15;
input 	A_mul_src1_16;
input 	A_mul_src1_17;
input 	A_mul_src1_18;
input 	A_mul_src1_19;
input 	A_mul_src1_20;
input 	A_mul_src1_21;
input 	A_mul_src1_22;
input 	A_mul_src1_23;
input 	A_mul_src1_24;
input 	A_mul_src1_25;
input 	A_mul_src1_26;
input 	A_mul_src1_27;
input 	A_mul_src1_28;
input 	A_mul_src1_29;
input 	A_mul_src1_30;
input 	A_mul_src1_31;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
output 	data_out_wire_2;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_0;
output 	data_out_wire_15;
output 	data_out_wire_14;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[21]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[20]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[25]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[17]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[24]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[16]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[27]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[19]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[26]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[18]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[23]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[22]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[29]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[30]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[31]~q ;
wire \the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ;
wire \the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[28]~q ;
wire \Add0~2 ;
wire \Add0~6 ;
wire \Add0~10 ;
wire \Add0~14 ;
wire \Add0~18 ;
wire \Add0~22 ;
wire \Add0~26 ;
wire \Add0~30 ;
wire \Add0~34 ;
wire \Add0~38 ;
wire \Add0~42 ;
wire \Add0~46 ;
wire \Add0~50 ;
wire \Add0~54 ;
wire \Add0~62 ;


embedded_system_altera_mult_add the_altmult_add_part_1(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_0(A_mul_src1_0),
	.A_mul_src1_1(A_mul_src1_1),
	.A_mul_src1_2(A_mul_src1_2),
	.A_mul_src1_3(A_mul_src1_3),
	.A_mul_src1_4(A_mul_src1_4),
	.A_mul_src1_5(A_mul_src1_5),
	.A_mul_src1_6(A_mul_src1_6),
	.A_mul_src1_7(A_mul_src1_7),
	.A_mul_src1_8(A_mul_src1_8),
	.A_mul_src1_9(A_mul_src1_9),
	.A_mul_src1_10(A_mul_src1_10),
	.A_mul_src1_11(A_mul_src1_11),
	.A_mul_src1_12(A_mul_src1_12),
	.A_mul_src1_13(A_mul_src1_13),
	.A_mul_src1_14(A_mul_src1_14),
	.A_mul_src1_15(A_mul_src1_15),
	.hq3myc14108phmpo7y7qmhbp98hy0vq(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_21(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[21]~q ),
	.data_out_wire_20(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[20]~q ),
	.data_out_wire_25(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[25]~q ),
	.data_out_wire_17(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[17]~q ),
	.data_out_wire_24(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[24]~q ),
	.data_out_wire_16(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[16]~q ),
	.data_out_wire_27(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[27]~q ),
	.data_out_wire_19(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[19]~q ),
	.data_out_wire_26(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[26]~q ),
	.data_out_wire_18(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[18]~q ),
	.data_out_wire_23(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[23]~q ),
	.data_out_wire_22(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[22]~q ),
	.data_out_wire_29(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[29]~q ),
	.data_out_wire_30(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[30]~q ),
	.data_out_wire_31(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[31]~q ),
	.data_out_wire_28(\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[28]~q ),
	.clk_clk(clk_clk));

embedded_system_altera_mult_add_1 the_altmult_add_part_2(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_16(A_mul_src1_16),
	.A_mul_src1_17(A_mul_src1_17),
	.A_mul_src1_18(A_mul_src1_18),
	.A_mul_src1_19(A_mul_src1_19),
	.A_mul_src1_20(A_mul_src1_20),
	.A_mul_src1_21(A_mul_src1_21),
	.A_mul_src1_22(A_mul_src1_22),
	.A_mul_src1_23(A_mul_src1_23),
	.A_mul_src1_24(A_mul_src1_24),
	.A_mul_src1_25(A_mul_src1_25),
	.A_mul_src1_26(A_mul_src1_26),
	.A_mul_src1_27(A_mul_src1_27),
	.A_mul_src1_28(A_mul_src1_28),
	.A_mul_src1_29(A_mul_src1_29),
	.A_mul_src1_30(A_mul_src1_30),
	.A_mul_src1_31(A_mul_src1_31),
	.hq3myc14108phmpo7y7qmhbp98hy0vq(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.data_out_wire_5(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.data_out_wire_4(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.data_out_wire_9(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.data_out_wire_1(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.data_out_wire_8(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.data_out_wire_0(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.data_out_wire_11(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.data_out_wire_3(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.data_out_wire_10(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.data_out_wire_2(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.data_out_wire_7(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.data_out_wire_6(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.data_out_wire_13(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.data_out_wire_14(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.data_out_wire_15(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.data_out_wire_12(\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.clk_clk(clk_clk));

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[5]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[21]~q ),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add0),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[4]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[20]~q ),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add01),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[9]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[25]~q ),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add02),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[1]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[17]~q ),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add03),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[8]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[24]~q ),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add04),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[0]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[16]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Add05),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[11]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[27]~q ),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add06),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[3]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[19]~q ),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add07),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[10]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[26]~q ),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add08),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

cyclonev_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[2]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[18]~q ),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add09),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

cyclonev_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[7]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[23]~q ),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add010),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

cyclonev_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[6]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[22]~q ),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add011),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

cyclonev_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[13]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[29]~q ),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add012),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

cyclonev_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[14]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[30]~q ),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add013),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

cyclonev_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[15]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[31]~q ),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add014),
	.cout(),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

cyclonev_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\the_altmult_add_part_2|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[12]~q ),
	.datae(gnd),
	.dataf(!\the_altmult_add_part_1|auto_generated|altera_mult_add_rtl1|multiplier_block|multiplier_register_block_0|data_out_wire[28]~q ),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(Add015),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

endmodule

module embedded_system_altera_mult_add (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_0,
	A_mul_src1_1,
	A_mul_src1_2,
	A_mul_src1_3,
	A_mul_src1_4,
	A_mul_src1_5,
	A_mul_src1_6,
	A_mul_src1_7,
	A_mul_src1_8,
	A_mul_src1_9,
	A_mul_src1_10,
	A_mul_src1_11,
	A_mul_src1_12,
	A_mul_src1_13,
	A_mul_src1_14,
	A_mul_src1_15,
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	data_out_wire_2,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_0,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_21,
	data_out_wire_20,
	data_out_wire_25,
	data_out_wire_17,
	data_out_wire_24,
	data_out_wire_16,
	data_out_wire_27,
	data_out_wire_19,
	data_out_wire_26,
	data_out_wire_18,
	data_out_wire_23,
	data_out_wire_22,
	data_out_wire_29,
	data_out_wire_30,
	data_out_wire_31,
	data_out_wire_28,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_0;
input 	A_mul_src1_1;
input 	A_mul_src1_2;
input 	A_mul_src1_3;
input 	A_mul_src1_4;
input 	A_mul_src1_5;
input 	A_mul_src1_6;
input 	A_mul_src1_7;
input 	A_mul_src1_8;
input 	A_mul_src1_9;
input 	A_mul_src1_10;
input 	A_mul_src1_11;
input 	A_mul_src1_12;
input 	A_mul_src1_13;
input 	A_mul_src1_14;
input 	A_mul_src1_15;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
output 	data_out_wire_2;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_0;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_21;
output 	data_out_wire_20;
output 	data_out_wire_25;
output 	data_out_wire_17;
output 	data_out_wire_24;
output 	data_out_wire_16;
output 	data_out_wire_27;
output 	data_out_wire_19;
output 	data_out_wire_26;
output 	data_out_wire_18;
output 	data_out_wire_23;
output 	data_out_wire_22;
output 	data_out_wire_29;
output 	data_out_wire_30;
output 	data_out_wire_31;
output 	data_out_wire_28;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altera_mult_add_ujt2 auto_generated(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_0(A_mul_src1_0),
	.A_mul_src1_1(A_mul_src1_1),
	.A_mul_src1_2(A_mul_src1_2),
	.A_mul_src1_3(A_mul_src1_3),
	.A_mul_src1_4(A_mul_src1_4),
	.A_mul_src1_5(A_mul_src1_5),
	.A_mul_src1_6(A_mul_src1_6),
	.A_mul_src1_7(A_mul_src1_7),
	.A_mul_src1_8(A_mul_src1_8),
	.A_mul_src1_9(A_mul_src1_9),
	.A_mul_src1_10(A_mul_src1_10),
	.A_mul_src1_11(A_mul_src1_11),
	.A_mul_src1_12(A_mul_src1_12),
	.A_mul_src1_13(A_mul_src1_13),
	.A_mul_src1_14(A_mul_src1_14),
	.A_mul_src1_15(A_mul_src1_15),
	.hq3myc14108phmpo7y7qmhbp98hy0vq(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_29(data_out_wire_29),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_31(data_out_wire_31),
	.data_out_wire_28(data_out_wire_28),
	.clk_clk(clk_clk));

endmodule

module embedded_system_altera_mult_add_ujt2 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_0,
	A_mul_src1_1,
	A_mul_src1_2,
	A_mul_src1_3,
	A_mul_src1_4,
	A_mul_src1_5,
	A_mul_src1_6,
	A_mul_src1_7,
	A_mul_src1_8,
	A_mul_src1_9,
	A_mul_src1_10,
	A_mul_src1_11,
	A_mul_src1_12,
	A_mul_src1_13,
	A_mul_src1_14,
	A_mul_src1_15,
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	data_out_wire_2,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_0,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_21,
	data_out_wire_20,
	data_out_wire_25,
	data_out_wire_17,
	data_out_wire_24,
	data_out_wire_16,
	data_out_wire_27,
	data_out_wire_19,
	data_out_wire_26,
	data_out_wire_18,
	data_out_wire_23,
	data_out_wire_22,
	data_out_wire_29,
	data_out_wire_30,
	data_out_wire_31,
	data_out_wire_28,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_0;
input 	A_mul_src1_1;
input 	A_mul_src1_2;
input 	A_mul_src1_3;
input 	A_mul_src1_4;
input 	A_mul_src1_5;
input 	A_mul_src1_6;
input 	A_mul_src1_7;
input 	A_mul_src1_8;
input 	A_mul_src1_9;
input 	A_mul_src1_10;
input 	A_mul_src1_11;
input 	A_mul_src1_12;
input 	A_mul_src1_13;
input 	A_mul_src1_14;
input 	A_mul_src1_15;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
output 	data_out_wire_2;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_0;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_21;
output 	data_out_wire_20;
output 	data_out_wire_25;
output 	data_out_wire_17;
output 	data_out_wire_24;
output 	data_out_wire_16;
output 	data_out_wire_27;
output 	data_out_wire_19;
output 	data_out_wire_26;
output 	data_out_wire_18;
output 	data_out_wire_23;
output 	data_out_wire_22;
output 	data_out_wire_29;
output 	data_out_wire_30;
output 	data_out_wire_31;
output 	data_out_wire_28;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altera_mult_add_rtl_1 altera_mult_add_rtl1(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_0(A_mul_src1_0),
	.A_mul_src1_1(A_mul_src1_1),
	.A_mul_src1_2(A_mul_src1_2),
	.A_mul_src1_3(A_mul_src1_3),
	.A_mul_src1_4(A_mul_src1_4),
	.A_mul_src1_5(A_mul_src1_5),
	.A_mul_src1_6(A_mul_src1_6),
	.A_mul_src1_7(A_mul_src1_7),
	.A_mul_src1_8(A_mul_src1_8),
	.A_mul_src1_9(A_mul_src1_9),
	.A_mul_src1_10(A_mul_src1_10),
	.A_mul_src1_11(A_mul_src1_11),
	.A_mul_src1_12(A_mul_src1_12),
	.A_mul_src1_13(A_mul_src1_13),
	.A_mul_src1_14(A_mul_src1_14),
	.A_mul_src1_15(A_mul_src1_15),
	.hq3myc14108phmpo7y7qmhbp98hy0vq(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_29(data_out_wire_29),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_31(data_out_wire_31),
	.data_out_wire_28(data_out_wire_28),
	.clk_clk(clk_clk));

endmodule

module embedded_system_altera_mult_add_rtl_1 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_0,
	A_mul_src1_1,
	A_mul_src1_2,
	A_mul_src1_3,
	A_mul_src1_4,
	A_mul_src1_5,
	A_mul_src1_6,
	A_mul_src1_7,
	A_mul_src1_8,
	A_mul_src1_9,
	A_mul_src1_10,
	A_mul_src1_11,
	A_mul_src1_12,
	A_mul_src1_13,
	A_mul_src1_14,
	A_mul_src1_15,
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	data_out_wire_2,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_0,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_21,
	data_out_wire_20,
	data_out_wire_25,
	data_out_wire_17,
	data_out_wire_24,
	data_out_wire_16,
	data_out_wire_27,
	data_out_wire_19,
	data_out_wire_26,
	data_out_wire_18,
	data_out_wire_23,
	data_out_wire_22,
	data_out_wire_29,
	data_out_wire_30,
	data_out_wire_31,
	data_out_wire_28,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_0;
input 	A_mul_src1_1;
input 	A_mul_src1_2;
input 	A_mul_src1_3;
input 	A_mul_src1_4;
input 	A_mul_src1_5;
input 	A_mul_src1_6;
input 	A_mul_src1_7;
input 	A_mul_src1_8;
input 	A_mul_src1_9;
input 	A_mul_src1_10;
input 	A_mul_src1_11;
input 	A_mul_src1_12;
input 	A_mul_src1_13;
input 	A_mul_src1_14;
input 	A_mul_src1_15;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
output 	data_out_wire_2;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_0;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_21;
output 	data_out_wire_20;
output 	data_out_wire_25;
output 	data_out_wire_17;
output 	data_out_wire_24;
output 	data_out_wire_16;
output 	data_out_wire_27;
output 	data_out_wire_19;
output 	data_out_wire_26;
output 	data_out_wire_18;
output 	data_out_wire_23;
output 	data_out_wire_22;
output 	data_out_wire_29;
output 	data_out_wire_30;
output 	data_out_wire_31;
output 	data_out_wire_28;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_ama_multiplier_function multiplier_block(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_0(A_mul_src1_0),
	.A_mul_src1_1(A_mul_src1_1),
	.A_mul_src1_2(A_mul_src1_2),
	.A_mul_src1_3(A_mul_src1_3),
	.A_mul_src1_4(A_mul_src1_4),
	.A_mul_src1_5(A_mul_src1_5),
	.A_mul_src1_6(A_mul_src1_6),
	.A_mul_src1_7(A_mul_src1_7),
	.A_mul_src1_8(A_mul_src1_8),
	.A_mul_src1_9(A_mul_src1_9),
	.A_mul_src1_10(A_mul_src1_10),
	.A_mul_src1_11(A_mul_src1_11),
	.A_mul_src1_12(A_mul_src1_12),
	.A_mul_src1_13(A_mul_src1_13),
	.A_mul_src1_14(A_mul_src1_14),
	.A_mul_src1_15(A_mul_src1_15),
	.hq3myc14108phmpo7y7qmhbp98hy0vq(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_29(data_out_wire_29),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_31(data_out_wire_31),
	.data_out_wire_28(data_out_wire_28),
	.clk_clk(clk_clk));

endmodule

module embedded_system_ama_multiplier_function (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_0,
	A_mul_src1_1,
	A_mul_src1_2,
	A_mul_src1_3,
	A_mul_src1_4,
	A_mul_src1_5,
	A_mul_src1_6,
	A_mul_src1_7,
	A_mul_src1_8,
	A_mul_src1_9,
	A_mul_src1_10,
	A_mul_src1_11,
	A_mul_src1_12,
	A_mul_src1_13,
	A_mul_src1_14,
	A_mul_src1_15,
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	data_out_wire_2,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_0,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_21,
	data_out_wire_20,
	data_out_wire_25,
	data_out_wire_17,
	data_out_wire_24,
	data_out_wire_16,
	data_out_wire_27,
	data_out_wire_19,
	data_out_wire_26,
	data_out_wire_18,
	data_out_wire_23,
	data_out_wire_22,
	data_out_wire_29,
	data_out_wire_30,
	data_out_wire_31,
	data_out_wire_28,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_0;
input 	A_mul_src1_1;
input 	A_mul_src1_2;
input 	A_mul_src1_3;
input 	A_mul_src1_4;
input 	A_mul_src1_5;
input 	A_mul_src1_6;
input 	A_mul_src1_7;
input 	A_mul_src1_8;
input 	A_mul_src1_9;
input 	A_mul_src1_10;
input 	A_mul_src1_11;
input 	A_mul_src1_12;
input 	A_mul_src1_13;
input 	A_mul_src1_14;
input 	A_mul_src1_15;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
output 	data_out_wire_2;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_0;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_21;
output 	data_out_wire_20;
output 	data_out_wire_25;
output 	data_out_wire_17;
output 	data_out_wire_24;
output 	data_out_wire_16;
output 	data_out_wire_27;
output 	data_out_wire_19;
output 	data_out_wire_26;
output 	data_out_wire_18;
output 	data_out_wire_23;
output 	data_out_wire_22;
output 	data_out_wire_29;
output 	data_out_wire_30;
output 	data_out_wire_31;
output 	data_out_wire_28;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out_wire_0[0] ;
wire \data_out_wire_0[1] ;
wire \data_out_wire_0[2] ;
wire \data_out_wire_0[3] ;
wire \data_out_wire_0[4] ;
wire \data_out_wire_0[5] ;
wire \data_out_wire_0[6] ;
wire \data_out_wire_0[7] ;
wire \data_out_wire_0[8] ;
wire \data_out_wire_0[9] ;
wire \data_out_wire_0[10] ;
wire \data_out_wire_0[11] ;
wire \data_out_wire_0[12] ;
wire \data_out_wire_0[13] ;
wire \data_out_wire_0[14] ;
wire \data_out_wire_0[15] ;
wire \data_out_wire_0[16] ;
wire \data_out_wire_0[17] ;
wire \data_out_wire_0[18] ;
wire \data_out_wire_0[19] ;
wire \data_out_wire_0[20] ;
wire \data_out_wire_0[21] ;
wire \data_out_wire_0[22] ;
wire \data_out_wire_0[23] ;
wire \data_out_wire_0[24] ;
wire \data_out_wire_0[25] ;
wire \data_out_wire_0[26] ;
wire \data_out_wire_0[27] ;
wire \data_out_wire_0[28] ;
wire \data_out_wire_0[29] ;
wire \data_out_wire_0[30] ;
wire \data_out_wire_0[31] ;
wire \Mult0~8 ;
wire \Mult0~9 ;
wire \Mult0~10 ;
wire \Mult0~11 ;
wire \Mult0~12 ;
wire \Mult0~13 ;
wire \Mult0~14 ;
wire \Mult0~15 ;
wire \Mult0~16 ;
wire \Mult0~17 ;
wire \Mult0~18 ;
wire \Mult0~19 ;
wire \Mult0~20 ;
wire \Mult0~21 ;
wire \Mult0~22 ;
wire \Mult0~23 ;
wire \Mult0~24 ;
wire \Mult0~25 ;
wire \Mult0~26 ;
wire \Mult0~27 ;
wire \Mult0~28 ;
wire \Mult0~29 ;
wire \Mult0~30 ;
wire \Mult0~31 ;
wire \Mult0~32 ;
wire \Mult0~33 ;
wire \Mult0~34 ;
wire \Mult0~35 ;
wire \Mult0~36 ;
wire \Mult0~37 ;
wire \Mult0~38 ;
wire \Mult0~39 ;

wire [63:0] \Mult0~mac_RESULTA_bus ;

assign \data_out_wire_0[0]  = \Mult0~mac_RESULTA_bus [0];
assign \data_out_wire_0[1]  = \Mult0~mac_RESULTA_bus [1];
assign \data_out_wire_0[2]  = \Mult0~mac_RESULTA_bus [2];
assign \data_out_wire_0[3]  = \Mult0~mac_RESULTA_bus [3];
assign \data_out_wire_0[4]  = \Mult0~mac_RESULTA_bus [4];
assign \data_out_wire_0[5]  = \Mult0~mac_RESULTA_bus [5];
assign \data_out_wire_0[6]  = \Mult0~mac_RESULTA_bus [6];
assign \data_out_wire_0[7]  = \Mult0~mac_RESULTA_bus [7];
assign \data_out_wire_0[8]  = \Mult0~mac_RESULTA_bus [8];
assign \data_out_wire_0[9]  = \Mult0~mac_RESULTA_bus [9];
assign \data_out_wire_0[10]  = \Mult0~mac_RESULTA_bus [10];
assign \data_out_wire_0[11]  = \Mult0~mac_RESULTA_bus [11];
assign \data_out_wire_0[12]  = \Mult0~mac_RESULTA_bus [12];
assign \data_out_wire_0[13]  = \Mult0~mac_RESULTA_bus [13];
assign \data_out_wire_0[14]  = \Mult0~mac_RESULTA_bus [14];
assign \data_out_wire_0[15]  = \Mult0~mac_RESULTA_bus [15];
assign \data_out_wire_0[16]  = \Mult0~mac_RESULTA_bus [16];
assign \data_out_wire_0[17]  = \Mult0~mac_RESULTA_bus [17];
assign \data_out_wire_0[18]  = \Mult0~mac_RESULTA_bus [18];
assign \data_out_wire_0[19]  = \Mult0~mac_RESULTA_bus [19];
assign \data_out_wire_0[20]  = \Mult0~mac_RESULTA_bus [20];
assign \data_out_wire_0[21]  = \Mult0~mac_RESULTA_bus [21];
assign \data_out_wire_0[22]  = \Mult0~mac_RESULTA_bus [22];
assign \data_out_wire_0[23]  = \Mult0~mac_RESULTA_bus [23];
assign \data_out_wire_0[24]  = \Mult0~mac_RESULTA_bus [24];
assign \data_out_wire_0[25]  = \Mult0~mac_RESULTA_bus [25];
assign \data_out_wire_0[26]  = \Mult0~mac_RESULTA_bus [26];
assign \data_out_wire_0[27]  = \Mult0~mac_RESULTA_bus [27];
assign \data_out_wire_0[28]  = \Mult0~mac_RESULTA_bus [28];
assign \data_out_wire_0[29]  = \Mult0~mac_RESULTA_bus [29];
assign \data_out_wire_0[30]  = \Mult0~mac_RESULTA_bus [30];
assign \data_out_wire_0[31]  = \Mult0~mac_RESULTA_bus [31];
assign \Mult0~8  = \Mult0~mac_RESULTA_bus [32];
assign \Mult0~9  = \Mult0~mac_RESULTA_bus [33];
assign \Mult0~10  = \Mult0~mac_RESULTA_bus [34];
assign \Mult0~11  = \Mult0~mac_RESULTA_bus [35];
assign \Mult0~12  = \Mult0~mac_RESULTA_bus [36];
assign \Mult0~13  = \Mult0~mac_RESULTA_bus [37];
assign \Mult0~14  = \Mult0~mac_RESULTA_bus [38];
assign \Mult0~15  = \Mult0~mac_RESULTA_bus [39];
assign \Mult0~16  = \Mult0~mac_RESULTA_bus [40];
assign \Mult0~17  = \Mult0~mac_RESULTA_bus [41];
assign \Mult0~18  = \Mult0~mac_RESULTA_bus [42];
assign \Mult0~19  = \Mult0~mac_RESULTA_bus [43];
assign \Mult0~20  = \Mult0~mac_RESULTA_bus [44];
assign \Mult0~21  = \Mult0~mac_RESULTA_bus [45];
assign \Mult0~22  = \Mult0~mac_RESULTA_bus [46];
assign \Mult0~23  = \Mult0~mac_RESULTA_bus [47];
assign \Mult0~24  = \Mult0~mac_RESULTA_bus [48];
assign \Mult0~25  = \Mult0~mac_RESULTA_bus [49];
assign \Mult0~26  = \Mult0~mac_RESULTA_bus [50];
assign \Mult0~27  = \Mult0~mac_RESULTA_bus [51];
assign \Mult0~28  = \Mult0~mac_RESULTA_bus [52];
assign \Mult0~29  = \Mult0~mac_RESULTA_bus [53];
assign \Mult0~30  = \Mult0~mac_RESULTA_bus [54];
assign \Mult0~31  = \Mult0~mac_RESULTA_bus [55];
assign \Mult0~32  = \Mult0~mac_RESULTA_bus [56];
assign \Mult0~33  = \Mult0~mac_RESULTA_bus [57];
assign \Mult0~34  = \Mult0~mac_RESULTA_bus [58];
assign \Mult0~35  = \Mult0~mac_RESULTA_bus [59];
assign \Mult0~36  = \Mult0~mac_RESULTA_bus [60];
assign \Mult0~37  = \Mult0~mac_RESULTA_bus [61];
assign \Mult0~38  = \Mult0~mac_RESULTA_bus [62];
assign \Mult0~39  = \Mult0~mac_RESULTA_bus [63];

embedded_system_ama_register_function_12 multiplier_register_block_0(
	.data_in({gnd,gnd,\data_out_wire_0[31] ,\data_out_wire_0[30] ,\data_out_wire_0[29] ,\data_out_wire_0[28] ,\data_out_wire_0[27] ,\data_out_wire_0[26] ,\data_out_wire_0[25] ,\data_out_wire_0[24] ,\data_out_wire_0[23] ,\data_out_wire_0[22] ,\data_out_wire_0[21] ,
\data_out_wire_0[20] ,\data_out_wire_0[19] ,\data_out_wire_0[18] ,\data_out_wire_0[17] ,\data_out_wire_0[16] ,\data_out_wire_0[15] ,\data_out_wire_0[14] ,\data_out_wire_0[13] ,\data_out_wire_0[12] ,\data_out_wire_0[11] ,\data_out_wire_0[10] ,\data_out_wire_0[9] ,
\data_out_wire_0[8] ,\data_out_wire_0[7] ,\data_out_wire_0[6] ,\data_out_wire_0[5] ,\data_out_wire_0[4] ,\data_out_wire_0[3] ,\data_out_wire_0[2] ,\data_out_wire_0[1] ,\data_out_wire_0[0] }),
	.aclr({gnd,gnd,gnd,hq3myc14108phmpo7y7qmhbp98hy0vq}),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_12(data_out_wire_12),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_21(data_out_wire_21),
	.data_out_wire_20(data_out_wire_20),
	.data_out_wire_25(data_out_wire_25),
	.data_out_wire_17(data_out_wire_17),
	.data_out_wire_24(data_out_wire_24),
	.data_out_wire_16(data_out_wire_16),
	.data_out_wire_27(data_out_wire_27),
	.data_out_wire_19(data_out_wire_19),
	.data_out_wire_26(data_out_wire_26),
	.data_out_wire_18(data_out_wire_18),
	.data_out_wire_23(data_out_wire_23),
	.data_out_wire_22(data_out_wire_22),
	.data_out_wire_29(data_out_wire_29),
	.data_out_wire_30(data_out_wire_30),
	.data_out_wire_31(data_out_wire_31),
	.data_out_wire_28(data_out_wire_28),
	.clock({gnd,gnd,gnd,clk_clk}));

cyclonev_mac \Mult0~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_mul_src2_15,A_mul_src2_14,A_mul_src2_13,A_mul_src2_12,A_mul_src2_11,A_mul_src2_10,A_mul_src2_9,A_mul_src2_8,A_mul_src2_7,A_mul_src2_6,A_mul_src2_5,A_mul_src2_4,A_mul_src2_3,A_mul_src2_2,A_mul_src2_1,A_mul_src2_0}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_mul_src1_15,A_mul_src1_14,A_mul_src1_13,A_mul_src1_12,A_mul_src1_11,A_mul_src1_10,A_mul_src1_9,A_mul_src1_8,A_mul_src1_7,A_mul_src1_6,A_mul_src1_5,A_mul_src1_4,A_mul_src1_3,A_mul_src1_2,A_mul_src1_1,A_mul_src1_0}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Mult0~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Mult0~mac .accumulate_clock = "none";
defparam \Mult0~mac .ax_clock = "none";
defparam \Mult0~mac .ax_width = 16;
defparam \Mult0~mac .ay_scan_in_clock = "none";
defparam \Mult0~mac .ay_scan_in_width = 16;
defparam \Mult0~mac .ay_use_scan_in = "false";
defparam \Mult0~mac .az_clock = "none";
defparam \Mult0~mac .bx_clock = "none";
defparam \Mult0~mac .by_clock = "none";
defparam \Mult0~mac .by_use_scan_in = "false";
defparam \Mult0~mac .bz_clock = "none";
defparam \Mult0~mac .coef_a_0 = 0;
defparam \Mult0~mac .coef_a_1 = 0;
defparam \Mult0~mac .coef_a_2 = 0;
defparam \Mult0~mac .coef_a_3 = 0;
defparam \Mult0~mac .coef_a_4 = 0;
defparam \Mult0~mac .coef_a_5 = 0;
defparam \Mult0~mac .coef_a_6 = 0;
defparam \Mult0~mac .coef_a_7 = 0;
defparam \Mult0~mac .coef_b_0 = 0;
defparam \Mult0~mac .coef_b_1 = 0;
defparam \Mult0~mac .coef_b_2 = 0;
defparam \Mult0~mac .coef_b_3 = 0;
defparam \Mult0~mac .coef_b_4 = 0;
defparam \Mult0~mac .coef_b_5 = 0;
defparam \Mult0~mac .coef_b_6 = 0;
defparam \Mult0~mac .coef_b_7 = 0;
defparam \Mult0~mac .coef_sel_a_clock = "none";
defparam \Mult0~mac .coef_sel_b_clock = "none";
defparam \Mult0~mac .delay_scan_out_ay = "false";
defparam \Mult0~mac .delay_scan_out_by = "false";
defparam \Mult0~mac .enable_double_accum = "false";
defparam \Mult0~mac .load_const_clock = "none";
defparam \Mult0~mac .load_const_value = 0;
defparam \Mult0~mac .mode_sub_location = 0;
defparam \Mult0~mac .negate_clock = "none";
defparam \Mult0~mac .operand_source_max = "input";
defparam \Mult0~mac .operand_source_may = "input";
defparam \Mult0~mac .operand_source_mbx = "input";
defparam \Mult0~mac .operand_source_mby = "input";
defparam \Mult0~mac .operation_mode = "m18x18_full";
defparam \Mult0~mac .output_clock = "none";
defparam \Mult0~mac .preadder_subtract_a = "false";
defparam \Mult0~mac .preadder_subtract_b = "false";
defparam \Mult0~mac .result_a_width = 64;
defparam \Mult0~mac .signed_max = "false";
defparam \Mult0~mac .signed_may = "false";
defparam \Mult0~mac .signed_mbx = "false";
defparam \Mult0~mac .signed_mby = "false";
defparam \Mult0~mac .sub_clock = "none";
defparam \Mult0~mac .use_chainadder = "false";

endmodule

module embedded_system_ama_register_function_12 (
	data_in,
	aclr,
	data_out_wire_2,
	data_out_wire_13,
	data_out_wire_12,
	data_out_wire_11,
	data_out_wire_10,
	data_out_wire_9,
	data_out_wire_8,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_3,
	data_out_wire_1,
	data_out_wire_0,
	data_out_wire_15,
	data_out_wire_14,
	data_out_wire_21,
	data_out_wire_20,
	data_out_wire_25,
	data_out_wire_17,
	data_out_wire_24,
	data_out_wire_16,
	data_out_wire_27,
	data_out_wire_19,
	data_out_wire_26,
	data_out_wire_18,
	data_out_wire_23,
	data_out_wire_22,
	data_out_wire_29,
	data_out_wire_30,
	data_out_wire_31,
	data_out_wire_28,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[33:0] data_in;
input 	[3:0] aclr;
output 	data_out_wire_2;
output 	data_out_wire_13;
output 	data_out_wire_12;
output 	data_out_wire_11;
output 	data_out_wire_10;
output 	data_out_wire_9;
output 	data_out_wire_8;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_3;
output 	data_out_wire_1;
output 	data_out_wire_0;
output 	data_out_wire_15;
output 	data_out_wire_14;
output 	data_out_wire_21;
output 	data_out_wire_20;
output 	data_out_wire_25;
output 	data_out_wire_17;
output 	data_out_wire_24;
output 	data_out_wire_16;
output 	data_out_wire_27;
output 	data_out_wire_19;
output 	data_out_wire_26;
output 	data_out_wire_18;
output 	data_out_wire_23;
output 	data_out_wire_22;
output 	data_out_wire_29;
output 	data_out_wire_30;
output 	data_out_wire_31;
output 	data_out_wire_28;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \data_out_wire[2] (
	.clk(clock[0]),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_2),
	.prn(vcc));
defparam \data_out_wire[2] .is_wysiwyg = "true";
defparam \data_out_wire[2] .power_up = "low";

dffeas \data_out_wire[13] (
	.clk(clock[0]),
	.d(data_in[13]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_13),
	.prn(vcc));
defparam \data_out_wire[13] .is_wysiwyg = "true";
defparam \data_out_wire[13] .power_up = "low";

dffeas \data_out_wire[12] (
	.clk(clock[0]),
	.d(data_in[12]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_12),
	.prn(vcc));
defparam \data_out_wire[12] .is_wysiwyg = "true";
defparam \data_out_wire[12] .power_up = "low";

dffeas \data_out_wire[11] (
	.clk(clock[0]),
	.d(data_in[11]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_11),
	.prn(vcc));
defparam \data_out_wire[11] .is_wysiwyg = "true";
defparam \data_out_wire[11] .power_up = "low";

dffeas \data_out_wire[10] (
	.clk(clock[0]),
	.d(data_in[10]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_10),
	.prn(vcc));
defparam \data_out_wire[10] .is_wysiwyg = "true";
defparam \data_out_wire[10] .power_up = "low";

dffeas \data_out_wire[9] (
	.clk(clock[0]),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_9),
	.prn(vcc));
defparam \data_out_wire[9] .is_wysiwyg = "true";
defparam \data_out_wire[9] .power_up = "low";

dffeas \data_out_wire[8] (
	.clk(clock[0]),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_8),
	.prn(vcc));
defparam \data_out_wire[8] .is_wysiwyg = "true";
defparam \data_out_wire[8] .power_up = "low";

dffeas \data_out_wire[7] (
	.clk(clock[0]),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_7),
	.prn(vcc));
defparam \data_out_wire[7] .is_wysiwyg = "true";
defparam \data_out_wire[7] .power_up = "low";

dffeas \data_out_wire[6] (
	.clk(clock[0]),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_6),
	.prn(vcc));
defparam \data_out_wire[6] .is_wysiwyg = "true";
defparam \data_out_wire[6] .power_up = "low";

dffeas \data_out_wire[5] (
	.clk(clock[0]),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_5),
	.prn(vcc));
defparam \data_out_wire[5] .is_wysiwyg = "true";
defparam \data_out_wire[5] .power_up = "low";

dffeas \data_out_wire[4] (
	.clk(clock[0]),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_4),
	.prn(vcc));
defparam \data_out_wire[4] .is_wysiwyg = "true";
defparam \data_out_wire[4] .power_up = "low";

dffeas \data_out_wire[3] (
	.clk(clock[0]),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_3),
	.prn(vcc));
defparam \data_out_wire[3] .is_wysiwyg = "true";
defparam \data_out_wire[3] .power_up = "low";

dffeas \data_out_wire[1] (
	.clk(clock[0]),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_1),
	.prn(vcc));
defparam \data_out_wire[1] .is_wysiwyg = "true";
defparam \data_out_wire[1] .power_up = "low";

dffeas \data_out_wire[0] (
	.clk(clock[0]),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_0),
	.prn(vcc));
defparam \data_out_wire[0] .is_wysiwyg = "true";
defparam \data_out_wire[0] .power_up = "low";

dffeas \data_out_wire[15] (
	.clk(clock[0]),
	.d(data_in[15]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_15),
	.prn(vcc));
defparam \data_out_wire[15] .is_wysiwyg = "true";
defparam \data_out_wire[15] .power_up = "low";

dffeas \data_out_wire[14] (
	.clk(clock[0]),
	.d(data_in[14]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_14),
	.prn(vcc));
defparam \data_out_wire[14] .is_wysiwyg = "true";
defparam \data_out_wire[14] .power_up = "low";

dffeas \data_out_wire[21] (
	.clk(clock[0]),
	.d(data_in[21]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_21),
	.prn(vcc));
defparam \data_out_wire[21] .is_wysiwyg = "true";
defparam \data_out_wire[21] .power_up = "low";

dffeas \data_out_wire[20] (
	.clk(clock[0]),
	.d(data_in[20]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_20),
	.prn(vcc));
defparam \data_out_wire[20] .is_wysiwyg = "true";
defparam \data_out_wire[20] .power_up = "low";

dffeas \data_out_wire[25] (
	.clk(clock[0]),
	.d(data_in[25]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_25),
	.prn(vcc));
defparam \data_out_wire[25] .is_wysiwyg = "true";
defparam \data_out_wire[25] .power_up = "low";

dffeas \data_out_wire[17] (
	.clk(clock[0]),
	.d(data_in[17]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_17),
	.prn(vcc));
defparam \data_out_wire[17] .is_wysiwyg = "true";
defparam \data_out_wire[17] .power_up = "low";

dffeas \data_out_wire[24] (
	.clk(clock[0]),
	.d(data_in[24]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_24),
	.prn(vcc));
defparam \data_out_wire[24] .is_wysiwyg = "true";
defparam \data_out_wire[24] .power_up = "low";

dffeas \data_out_wire[16] (
	.clk(clock[0]),
	.d(data_in[16]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_16),
	.prn(vcc));
defparam \data_out_wire[16] .is_wysiwyg = "true";
defparam \data_out_wire[16] .power_up = "low";

dffeas \data_out_wire[27] (
	.clk(clock[0]),
	.d(data_in[27]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_27),
	.prn(vcc));
defparam \data_out_wire[27] .is_wysiwyg = "true";
defparam \data_out_wire[27] .power_up = "low";

dffeas \data_out_wire[19] (
	.clk(clock[0]),
	.d(data_in[19]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_19),
	.prn(vcc));
defparam \data_out_wire[19] .is_wysiwyg = "true";
defparam \data_out_wire[19] .power_up = "low";

dffeas \data_out_wire[26] (
	.clk(clock[0]),
	.d(data_in[26]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_26),
	.prn(vcc));
defparam \data_out_wire[26] .is_wysiwyg = "true";
defparam \data_out_wire[26] .power_up = "low";

dffeas \data_out_wire[18] (
	.clk(clock[0]),
	.d(data_in[18]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_18),
	.prn(vcc));
defparam \data_out_wire[18] .is_wysiwyg = "true";
defparam \data_out_wire[18] .power_up = "low";

dffeas \data_out_wire[23] (
	.clk(clock[0]),
	.d(data_in[23]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_23),
	.prn(vcc));
defparam \data_out_wire[23] .is_wysiwyg = "true";
defparam \data_out_wire[23] .power_up = "low";

dffeas \data_out_wire[22] (
	.clk(clock[0]),
	.d(data_in[22]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_22),
	.prn(vcc));
defparam \data_out_wire[22] .is_wysiwyg = "true";
defparam \data_out_wire[22] .power_up = "low";

dffeas \data_out_wire[29] (
	.clk(clock[0]),
	.d(data_in[29]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_29),
	.prn(vcc));
defparam \data_out_wire[29] .is_wysiwyg = "true";
defparam \data_out_wire[29] .power_up = "low";

dffeas \data_out_wire[30] (
	.clk(clock[0]),
	.d(data_in[30]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_30),
	.prn(vcc));
defparam \data_out_wire[30] .is_wysiwyg = "true";
defparam \data_out_wire[30] .power_up = "low";

dffeas \data_out_wire[31] (
	.clk(clock[0]),
	.d(data_in[31]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_31),
	.prn(vcc));
defparam \data_out_wire[31] .is_wysiwyg = "true";
defparam \data_out_wire[31] .power_up = "low";

dffeas \data_out_wire[28] (
	.clk(clock[0]),
	.d(data_in[28]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_28),
	.prn(vcc));
defparam \data_out_wire[28] .is_wysiwyg = "true";
defparam \data_out_wire[28] .power_up = "low";

endmodule

module embedded_system_altera_mult_add_1 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_16,
	A_mul_src1_17,
	A_mul_src1_18,
	A_mul_src1_19,
	A_mul_src1_20,
	A_mul_src1_21,
	A_mul_src1_22,
	A_mul_src1_23,
	A_mul_src1_24,
	A_mul_src1_25,
	A_mul_src1_26,
	A_mul_src1_27,
	A_mul_src1_28,
	A_mul_src1_29,
	A_mul_src1_30,
	A_mul_src1_31,
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_9,
	data_out_wire_1,
	data_out_wire_8,
	data_out_wire_0,
	data_out_wire_11,
	data_out_wire_3,
	data_out_wire_10,
	data_out_wire_2,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_15,
	data_out_wire_12,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_16;
input 	A_mul_src1_17;
input 	A_mul_src1_18;
input 	A_mul_src1_19;
input 	A_mul_src1_20;
input 	A_mul_src1_21;
input 	A_mul_src1_22;
input 	A_mul_src1_23;
input 	A_mul_src1_24;
input 	A_mul_src1_25;
input 	A_mul_src1_26;
input 	A_mul_src1_27;
input 	A_mul_src1_28;
input 	A_mul_src1_29;
input 	A_mul_src1_30;
input 	A_mul_src1_31;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_9;
output 	data_out_wire_1;
output 	data_out_wire_8;
output 	data_out_wire_0;
output 	data_out_wire_11;
output 	data_out_wire_3;
output 	data_out_wire_10;
output 	data_out_wire_2;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_15;
output 	data_out_wire_12;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altera_mult_add_0kt2 auto_generated(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_16(A_mul_src1_16),
	.A_mul_src1_17(A_mul_src1_17),
	.A_mul_src1_18(A_mul_src1_18),
	.A_mul_src1_19(A_mul_src1_19),
	.A_mul_src1_20(A_mul_src1_20),
	.A_mul_src1_21(A_mul_src1_21),
	.A_mul_src1_22(A_mul_src1_22),
	.A_mul_src1_23(A_mul_src1_23),
	.A_mul_src1_24(A_mul_src1_24),
	.A_mul_src1_25(A_mul_src1_25),
	.A_mul_src1_26(A_mul_src1_26),
	.A_mul_src1_27(A_mul_src1_27),
	.A_mul_src1_28(A_mul_src1_28),
	.A_mul_src1_29(A_mul_src1_29),
	.A_mul_src1_30(A_mul_src1_30),
	.A_mul_src1_31(A_mul_src1_31),
	.hq3myc14108phmpo7y7qmhbp98hy0vq(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_12(data_out_wire_12),
	.clk_clk(clk_clk));

endmodule

module embedded_system_altera_mult_add_0kt2 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_16,
	A_mul_src1_17,
	A_mul_src1_18,
	A_mul_src1_19,
	A_mul_src1_20,
	A_mul_src1_21,
	A_mul_src1_22,
	A_mul_src1_23,
	A_mul_src1_24,
	A_mul_src1_25,
	A_mul_src1_26,
	A_mul_src1_27,
	A_mul_src1_28,
	A_mul_src1_29,
	A_mul_src1_30,
	A_mul_src1_31,
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_9,
	data_out_wire_1,
	data_out_wire_8,
	data_out_wire_0,
	data_out_wire_11,
	data_out_wire_3,
	data_out_wire_10,
	data_out_wire_2,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_15,
	data_out_wire_12,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_16;
input 	A_mul_src1_17;
input 	A_mul_src1_18;
input 	A_mul_src1_19;
input 	A_mul_src1_20;
input 	A_mul_src1_21;
input 	A_mul_src1_22;
input 	A_mul_src1_23;
input 	A_mul_src1_24;
input 	A_mul_src1_25;
input 	A_mul_src1_26;
input 	A_mul_src1_27;
input 	A_mul_src1_28;
input 	A_mul_src1_29;
input 	A_mul_src1_30;
input 	A_mul_src1_31;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_9;
output 	data_out_wire_1;
output 	data_out_wire_8;
output 	data_out_wire_0;
output 	data_out_wire_11;
output 	data_out_wire_3;
output 	data_out_wire_10;
output 	data_out_wire_2;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_15;
output 	data_out_wire_12;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altera_mult_add_rtl_2 altera_mult_add_rtl1(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_16(A_mul_src1_16),
	.A_mul_src1_17(A_mul_src1_17),
	.A_mul_src1_18(A_mul_src1_18),
	.A_mul_src1_19(A_mul_src1_19),
	.A_mul_src1_20(A_mul_src1_20),
	.A_mul_src1_21(A_mul_src1_21),
	.A_mul_src1_22(A_mul_src1_22),
	.A_mul_src1_23(A_mul_src1_23),
	.A_mul_src1_24(A_mul_src1_24),
	.A_mul_src1_25(A_mul_src1_25),
	.A_mul_src1_26(A_mul_src1_26),
	.A_mul_src1_27(A_mul_src1_27),
	.A_mul_src1_28(A_mul_src1_28),
	.A_mul_src1_29(A_mul_src1_29),
	.A_mul_src1_30(A_mul_src1_30),
	.A_mul_src1_31(A_mul_src1_31),
	.hq3myc14108phmpo7y7qmhbp98hy0vq(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_12(data_out_wire_12),
	.clk_clk(clk_clk));

endmodule

module embedded_system_altera_mult_add_rtl_2 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_16,
	A_mul_src1_17,
	A_mul_src1_18,
	A_mul_src1_19,
	A_mul_src1_20,
	A_mul_src1_21,
	A_mul_src1_22,
	A_mul_src1_23,
	A_mul_src1_24,
	A_mul_src1_25,
	A_mul_src1_26,
	A_mul_src1_27,
	A_mul_src1_28,
	A_mul_src1_29,
	A_mul_src1_30,
	A_mul_src1_31,
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_9,
	data_out_wire_1,
	data_out_wire_8,
	data_out_wire_0,
	data_out_wire_11,
	data_out_wire_3,
	data_out_wire_10,
	data_out_wire_2,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_15,
	data_out_wire_12,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_16;
input 	A_mul_src1_17;
input 	A_mul_src1_18;
input 	A_mul_src1_19;
input 	A_mul_src1_20;
input 	A_mul_src1_21;
input 	A_mul_src1_22;
input 	A_mul_src1_23;
input 	A_mul_src1_24;
input 	A_mul_src1_25;
input 	A_mul_src1_26;
input 	A_mul_src1_27;
input 	A_mul_src1_28;
input 	A_mul_src1_29;
input 	A_mul_src1_30;
input 	A_mul_src1_31;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_9;
output 	data_out_wire_1;
output 	data_out_wire_8;
output 	data_out_wire_0;
output 	data_out_wire_11;
output 	data_out_wire_3;
output 	data_out_wire_10;
output 	data_out_wire_2;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_15;
output 	data_out_wire_12;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_ama_multiplier_function_1 multiplier_block(
	.A_mul_src2_0(A_mul_src2_0),
	.A_mul_src2_1(A_mul_src2_1),
	.A_mul_src2_2(A_mul_src2_2),
	.A_mul_src2_3(A_mul_src2_3),
	.A_mul_src2_4(A_mul_src2_4),
	.A_mul_src2_5(A_mul_src2_5),
	.A_mul_src2_6(A_mul_src2_6),
	.A_mul_src2_7(A_mul_src2_7),
	.A_mul_src2_8(A_mul_src2_8),
	.A_mul_src2_9(A_mul_src2_9),
	.A_mul_src2_10(A_mul_src2_10),
	.A_mul_src2_11(A_mul_src2_11),
	.A_mul_src2_12(A_mul_src2_12),
	.A_mul_src2_13(A_mul_src2_13),
	.A_mul_src2_14(A_mul_src2_14),
	.A_mul_src2_15(A_mul_src2_15),
	.A_mul_src1_16(A_mul_src1_16),
	.A_mul_src1_17(A_mul_src1_17),
	.A_mul_src1_18(A_mul_src1_18),
	.A_mul_src1_19(A_mul_src1_19),
	.A_mul_src1_20(A_mul_src1_20),
	.A_mul_src1_21(A_mul_src1_21),
	.A_mul_src1_22(A_mul_src1_22),
	.A_mul_src1_23(A_mul_src1_23),
	.A_mul_src1_24(A_mul_src1_24),
	.A_mul_src1_25(A_mul_src1_25),
	.A_mul_src1_26(A_mul_src1_26),
	.A_mul_src1_27(A_mul_src1_27),
	.A_mul_src1_28(A_mul_src1_28),
	.A_mul_src1_29(A_mul_src1_29),
	.A_mul_src1_30(A_mul_src1_30),
	.A_mul_src1_31(A_mul_src1_31),
	.hq3myc14108phmpo7y7qmhbp98hy0vq(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_12(data_out_wire_12),
	.clk_clk(clk_clk));

endmodule

module embedded_system_ama_multiplier_function_1 (
	A_mul_src2_0,
	A_mul_src2_1,
	A_mul_src2_2,
	A_mul_src2_3,
	A_mul_src2_4,
	A_mul_src2_5,
	A_mul_src2_6,
	A_mul_src2_7,
	A_mul_src2_8,
	A_mul_src2_9,
	A_mul_src2_10,
	A_mul_src2_11,
	A_mul_src2_12,
	A_mul_src2_13,
	A_mul_src2_14,
	A_mul_src2_15,
	A_mul_src1_16,
	A_mul_src1_17,
	A_mul_src1_18,
	A_mul_src1_19,
	A_mul_src1_20,
	A_mul_src1_21,
	A_mul_src1_22,
	A_mul_src1_23,
	A_mul_src1_24,
	A_mul_src1_25,
	A_mul_src1_26,
	A_mul_src1_27,
	A_mul_src1_28,
	A_mul_src1_29,
	A_mul_src1_30,
	A_mul_src1_31,
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_9,
	data_out_wire_1,
	data_out_wire_8,
	data_out_wire_0,
	data_out_wire_11,
	data_out_wire_3,
	data_out_wire_10,
	data_out_wire_2,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_15,
	data_out_wire_12,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	A_mul_src2_0;
input 	A_mul_src2_1;
input 	A_mul_src2_2;
input 	A_mul_src2_3;
input 	A_mul_src2_4;
input 	A_mul_src2_5;
input 	A_mul_src2_6;
input 	A_mul_src2_7;
input 	A_mul_src2_8;
input 	A_mul_src2_9;
input 	A_mul_src2_10;
input 	A_mul_src2_11;
input 	A_mul_src2_12;
input 	A_mul_src2_13;
input 	A_mul_src2_14;
input 	A_mul_src2_15;
input 	A_mul_src1_16;
input 	A_mul_src1_17;
input 	A_mul_src1_18;
input 	A_mul_src1_19;
input 	A_mul_src1_20;
input 	A_mul_src1_21;
input 	A_mul_src1_22;
input 	A_mul_src1_23;
input 	A_mul_src1_24;
input 	A_mul_src1_25;
input 	A_mul_src1_26;
input 	A_mul_src1_27;
input 	A_mul_src1_28;
input 	A_mul_src1_29;
input 	A_mul_src1_30;
input 	A_mul_src1_31;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_9;
output 	data_out_wire_1;
output 	data_out_wire_8;
output 	data_out_wire_0;
output 	data_out_wire_11;
output 	data_out_wire_3;
output 	data_out_wire_10;
output 	data_out_wire_2;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_15;
output 	data_out_wire_12;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \data_out_wire_0[0] ;
wire \data_out_wire_0[1] ;
wire \data_out_wire_0[2] ;
wire \data_out_wire_0[3] ;
wire \data_out_wire_0[4] ;
wire \data_out_wire_0[5] ;
wire \data_out_wire_0[6] ;
wire \data_out_wire_0[7] ;
wire \data_out_wire_0[8] ;
wire \data_out_wire_0[9] ;
wire \data_out_wire_0[10] ;
wire \data_out_wire_0[11] ;
wire \data_out_wire_0[12] ;
wire \data_out_wire_0[13] ;
wire \data_out_wire_0[14] ;
wire \data_out_wire_0[15] ;
wire \Mult0~8 ;
wire \Mult0~9 ;
wire \Mult0~10 ;
wire \Mult0~11 ;
wire \Mult0~12 ;
wire \Mult0~13 ;
wire \Mult0~14 ;
wire \Mult0~15 ;
wire \Mult0~16 ;
wire \Mult0~17 ;
wire \Mult0~18 ;
wire \Mult0~19 ;
wire \Mult0~20 ;
wire \Mult0~21 ;
wire \Mult0~22 ;
wire \Mult0~23 ;
wire \Mult0~24 ;
wire \Mult0~25 ;
wire \Mult0~26 ;
wire \Mult0~27 ;
wire \Mult0~28 ;
wire \Mult0~29 ;
wire \Mult0~30 ;
wire \Mult0~31 ;
wire \Mult0~32 ;
wire \Mult0~33 ;
wire \Mult0~34 ;
wire \Mult0~35 ;
wire \Mult0~36 ;
wire \Mult0~37 ;
wire \Mult0~38 ;
wire \Mult0~39 ;
wire \Mult0~40 ;
wire \Mult0~41 ;
wire \Mult0~42 ;
wire \Mult0~43 ;
wire \Mult0~44 ;
wire \Mult0~45 ;
wire \Mult0~46 ;
wire \Mult0~47 ;
wire \Mult0~48 ;
wire \Mult0~49 ;
wire \Mult0~50 ;
wire \Mult0~51 ;
wire \Mult0~52 ;
wire \Mult0~53 ;
wire \Mult0~54 ;
wire \Mult0~55 ;

wire [63:0] \Mult0~mac_RESULTA_bus ;

assign \data_out_wire_0[0]  = \Mult0~mac_RESULTA_bus [0];
assign \data_out_wire_0[1]  = \Mult0~mac_RESULTA_bus [1];
assign \data_out_wire_0[2]  = \Mult0~mac_RESULTA_bus [2];
assign \data_out_wire_0[3]  = \Mult0~mac_RESULTA_bus [3];
assign \data_out_wire_0[4]  = \Mult0~mac_RESULTA_bus [4];
assign \data_out_wire_0[5]  = \Mult0~mac_RESULTA_bus [5];
assign \data_out_wire_0[6]  = \Mult0~mac_RESULTA_bus [6];
assign \data_out_wire_0[7]  = \Mult0~mac_RESULTA_bus [7];
assign \data_out_wire_0[8]  = \Mult0~mac_RESULTA_bus [8];
assign \data_out_wire_0[9]  = \Mult0~mac_RESULTA_bus [9];
assign \data_out_wire_0[10]  = \Mult0~mac_RESULTA_bus [10];
assign \data_out_wire_0[11]  = \Mult0~mac_RESULTA_bus [11];
assign \data_out_wire_0[12]  = \Mult0~mac_RESULTA_bus [12];
assign \data_out_wire_0[13]  = \Mult0~mac_RESULTA_bus [13];
assign \data_out_wire_0[14]  = \Mult0~mac_RESULTA_bus [14];
assign \data_out_wire_0[15]  = \Mult0~mac_RESULTA_bus [15];
assign \Mult0~8  = \Mult0~mac_RESULTA_bus [16];
assign \Mult0~9  = \Mult0~mac_RESULTA_bus [17];
assign \Mult0~10  = \Mult0~mac_RESULTA_bus [18];
assign \Mult0~11  = \Mult0~mac_RESULTA_bus [19];
assign \Mult0~12  = \Mult0~mac_RESULTA_bus [20];
assign \Mult0~13  = \Mult0~mac_RESULTA_bus [21];
assign \Mult0~14  = \Mult0~mac_RESULTA_bus [22];
assign \Mult0~15  = \Mult0~mac_RESULTA_bus [23];
assign \Mult0~16  = \Mult0~mac_RESULTA_bus [24];
assign \Mult0~17  = \Mult0~mac_RESULTA_bus [25];
assign \Mult0~18  = \Mult0~mac_RESULTA_bus [26];
assign \Mult0~19  = \Mult0~mac_RESULTA_bus [27];
assign \Mult0~20  = \Mult0~mac_RESULTA_bus [28];
assign \Mult0~21  = \Mult0~mac_RESULTA_bus [29];
assign \Mult0~22  = \Mult0~mac_RESULTA_bus [30];
assign \Mult0~23  = \Mult0~mac_RESULTA_bus [31];
assign \Mult0~24  = \Mult0~mac_RESULTA_bus [32];
assign \Mult0~25  = \Mult0~mac_RESULTA_bus [33];
assign \Mult0~26  = \Mult0~mac_RESULTA_bus [34];
assign \Mult0~27  = \Mult0~mac_RESULTA_bus [35];
assign \Mult0~28  = \Mult0~mac_RESULTA_bus [36];
assign \Mult0~29  = \Mult0~mac_RESULTA_bus [37];
assign \Mult0~30  = \Mult0~mac_RESULTA_bus [38];
assign \Mult0~31  = \Mult0~mac_RESULTA_bus [39];
assign \Mult0~32  = \Mult0~mac_RESULTA_bus [40];
assign \Mult0~33  = \Mult0~mac_RESULTA_bus [41];
assign \Mult0~34  = \Mult0~mac_RESULTA_bus [42];
assign \Mult0~35  = \Mult0~mac_RESULTA_bus [43];
assign \Mult0~36  = \Mult0~mac_RESULTA_bus [44];
assign \Mult0~37  = \Mult0~mac_RESULTA_bus [45];
assign \Mult0~38  = \Mult0~mac_RESULTA_bus [46];
assign \Mult0~39  = \Mult0~mac_RESULTA_bus [47];
assign \Mult0~40  = \Mult0~mac_RESULTA_bus [48];
assign \Mult0~41  = \Mult0~mac_RESULTA_bus [49];
assign \Mult0~42  = \Mult0~mac_RESULTA_bus [50];
assign \Mult0~43  = \Mult0~mac_RESULTA_bus [51];
assign \Mult0~44  = \Mult0~mac_RESULTA_bus [52];
assign \Mult0~45  = \Mult0~mac_RESULTA_bus [53];
assign \Mult0~46  = \Mult0~mac_RESULTA_bus [54];
assign \Mult0~47  = \Mult0~mac_RESULTA_bus [55];
assign \Mult0~48  = \Mult0~mac_RESULTA_bus [56];
assign \Mult0~49  = \Mult0~mac_RESULTA_bus [57];
assign \Mult0~50  = \Mult0~mac_RESULTA_bus [58];
assign \Mult0~51  = \Mult0~mac_RESULTA_bus [59];
assign \Mult0~52  = \Mult0~mac_RESULTA_bus [60];
assign \Mult0~53  = \Mult0~mac_RESULTA_bus [61];
assign \Mult0~54  = \Mult0~mac_RESULTA_bus [62];
assign \Mult0~55  = \Mult0~mac_RESULTA_bus [63];

embedded_system_ama_register_function_31 multiplier_register_block_0(
	.data_in({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\data_out_wire_0[15] ,\data_out_wire_0[14] ,\data_out_wire_0[13] ,\data_out_wire_0[12] ,\data_out_wire_0[11] ,\data_out_wire_0[10] ,\data_out_wire_0[9] ,\data_out_wire_0[8] ,\data_out_wire_0[7] ,
\data_out_wire_0[6] ,\data_out_wire_0[5] ,\data_out_wire_0[4] ,\data_out_wire_0[3] ,\data_out_wire_0[2] ,\data_out_wire_0[1] ,\data_out_wire_0[0] }),
	.aclr({gnd,gnd,gnd,hq3myc14108phmpo7y7qmhbp98hy0vq}),
	.data_out_wire_5(data_out_wire_5),
	.data_out_wire_4(data_out_wire_4),
	.data_out_wire_9(data_out_wire_9),
	.data_out_wire_1(data_out_wire_1),
	.data_out_wire_8(data_out_wire_8),
	.data_out_wire_0(data_out_wire_0),
	.data_out_wire_11(data_out_wire_11),
	.data_out_wire_3(data_out_wire_3),
	.data_out_wire_10(data_out_wire_10),
	.data_out_wire_2(data_out_wire_2),
	.data_out_wire_7(data_out_wire_7),
	.data_out_wire_6(data_out_wire_6),
	.data_out_wire_13(data_out_wire_13),
	.data_out_wire_14(data_out_wire_14),
	.data_out_wire_15(data_out_wire_15),
	.data_out_wire_12(data_out_wire_12),
	.clock({gnd,gnd,gnd,clk_clk}));

cyclonev_mac \Mult0~mac (
	.sub(gnd),
	.negate(gnd),
	.accumulate(gnd),
	.loadconst(gnd),
	.ax({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_mul_src2_15,A_mul_src2_14,A_mul_src2_13,A_mul_src2_12,A_mul_src2_11,A_mul_src2_10,A_mul_src2_9,A_mul_src2_8,A_mul_src2_7,A_mul_src2_6,A_mul_src2_5,A_mul_src2_4,A_mul_src2_3,A_mul_src2_2,A_mul_src2_1,A_mul_src2_0}),
	.ay({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,A_mul_src1_31,A_mul_src1_30,A_mul_src1_29,A_mul_src1_28,A_mul_src1_27,A_mul_src1_26,A_mul_src1_25,A_mul_src1_24,A_mul_src1_23,A_mul_src1_22,A_mul_src1_21,A_mul_src1_20,A_mul_src1_19,A_mul_src1_18,A_mul_src1_17,A_mul_src1_16}),
	.az(26'b00000000000000000000000000),
	.bx(18'b000000000000000000),
	.by(19'b0000000000000000000),
	.bz(18'b000000000000000000),
	.coefsela(3'b000),
	.coefselb(3'b000),
	.clk(3'b000),
	.aclr(2'b00),
	.ena(3'b111),
	.scanin(27'b000000000000000000000000000),
	.chainin(1'b0),
	.dftout(),
	.resulta(\Mult0~mac_RESULTA_bus ),
	.resultb(),
	.scanout(),
	.chainout());
defparam \Mult0~mac .accumulate_clock = "none";
defparam \Mult0~mac .ax_clock = "none";
defparam \Mult0~mac .ax_width = 16;
defparam \Mult0~mac .ay_scan_in_clock = "none";
defparam \Mult0~mac .ay_scan_in_width = 16;
defparam \Mult0~mac .ay_use_scan_in = "false";
defparam \Mult0~mac .az_clock = "none";
defparam \Mult0~mac .bx_clock = "none";
defparam \Mult0~mac .by_clock = "none";
defparam \Mult0~mac .by_use_scan_in = "false";
defparam \Mult0~mac .bz_clock = "none";
defparam \Mult0~mac .coef_a_0 = 0;
defparam \Mult0~mac .coef_a_1 = 0;
defparam \Mult0~mac .coef_a_2 = 0;
defparam \Mult0~mac .coef_a_3 = 0;
defparam \Mult0~mac .coef_a_4 = 0;
defparam \Mult0~mac .coef_a_5 = 0;
defparam \Mult0~mac .coef_a_6 = 0;
defparam \Mult0~mac .coef_a_7 = 0;
defparam \Mult0~mac .coef_b_0 = 0;
defparam \Mult0~mac .coef_b_1 = 0;
defparam \Mult0~mac .coef_b_2 = 0;
defparam \Mult0~mac .coef_b_3 = 0;
defparam \Mult0~mac .coef_b_4 = 0;
defparam \Mult0~mac .coef_b_5 = 0;
defparam \Mult0~mac .coef_b_6 = 0;
defparam \Mult0~mac .coef_b_7 = 0;
defparam \Mult0~mac .coef_sel_a_clock = "none";
defparam \Mult0~mac .coef_sel_b_clock = "none";
defparam \Mult0~mac .delay_scan_out_ay = "false";
defparam \Mult0~mac .delay_scan_out_by = "false";
defparam \Mult0~mac .enable_double_accum = "false";
defparam \Mult0~mac .load_const_clock = "none";
defparam \Mult0~mac .load_const_value = 0;
defparam \Mult0~mac .mode_sub_location = 0;
defparam \Mult0~mac .negate_clock = "none";
defparam \Mult0~mac .operand_source_max = "input";
defparam \Mult0~mac .operand_source_may = "input";
defparam \Mult0~mac .operand_source_mbx = "input";
defparam \Mult0~mac .operand_source_mby = "input";
defparam \Mult0~mac .operation_mode = "m18x18_full";
defparam \Mult0~mac .output_clock = "none";
defparam \Mult0~mac .preadder_subtract_a = "false";
defparam \Mult0~mac .preadder_subtract_b = "false";
defparam \Mult0~mac .result_a_width = 64;
defparam \Mult0~mac .signed_max = "false";
defparam \Mult0~mac .signed_may = "false";
defparam \Mult0~mac .signed_mbx = "false";
defparam \Mult0~mac .signed_mby = "false";
defparam \Mult0~mac .sub_clock = "none";
defparam \Mult0~mac .use_chainadder = "false";

endmodule

module embedded_system_ama_register_function_31 (
	data_in,
	aclr,
	data_out_wire_5,
	data_out_wire_4,
	data_out_wire_9,
	data_out_wire_1,
	data_out_wire_8,
	data_out_wire_0,
	data_out_wire_11,
	data_out_wire_3,
	data_out_wire_10,
	data_out_wire_2,
	data_out_wire_7,
	data_out_wire_6,
	data_out_wire_13,
	data_out_wire_14,
	data_out_wire_15,
	data_out_wire_12,
	clock)/* synthesis synthesis_greybox=1 */;
input 	[33:0] data_in;
input 	[3:0] aclr;
output 	data_out_wire_5;
output 	data_out_wire_4;
output 	data_out_wire_9;
output 	data_out_wire_1;
output 	data_out_wire_8;
output 	data_out_wire_0;
output 	data_out_wire_11;
output 	data_out_wire_3;
output 	data_out_wire_10;
output 	data_out_wire_2;
output 	data_out_wire_7;
output 	data_out_wire_6;
output 	data_out_wire_13;
output 	data_out_wire_14;
output 	data_out_wire_15;
output 	data_out_wire_12;
input 	[3:0] clock;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \data_out_wire[5] (
	.clk(clock[0]),
	.d(data_in[5]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_5),
	.prn(vcc));
defparam \data_out_wire[5] .is_wysiwyg = "true";
defparam \data_out_wire[5] .power_up = "low";

dffeas \data_out_wire[4] (
	.clk(clock[0]),
	.d(data_in[4]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_4),
	.prn(vcc));
defparam \data_out_wire[4] .is_wysiwyg = "true";
defparam \data_out_wire[4] .power_up = "low";

dffeas \data_out_wire[9] (
	.clk(clock[0]),
	.d(data_in[9]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_9),
	.prn(vcc));
defparam \data_out_wire[9] .is_wysiwyg = "true";
defparam \data_out_wire[9] .power_up = "low";

dffeas \data_out_wire[1] (
	.clk(clock[0]),
	.d(data_in[1]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_1),
	.prn(vcc));
defparam \data_out_wire[1] .is_wysiwyg = "true";
defparam \data_out_wire[1] .power_up = "low";

dffeas \data_out_wire[8] (
	.clk(clock[0]),
	.d(data_in[8]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_8),
	.prn(vcc));
defparam \data_out_wire[8] .is_wysiwyg = "true";
defparam \data_out_wire[8] .power_up = "low";

dffeas \data_out_wire[0] (
	.clk(clock[0]),
	.d(data_in[0]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_0),
	.prn(vcc));
defparam \data_out_wire[0] .is_wysiwyg = "true";
defparam \data_out_wire[0] .power_up = "low";

dffeas \data_out_wire[11] (
	.clk(clock[0]),
	.d(data_in[11]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_11),
	.prn(vcc));
defparam \data_out_wire[11] .is_wysiwyg = "true";
defparam \data_out_wire[11] .power_up = "low";

dffeas \data_out_wire[3] (
	.clk(clock[0]),
	.d(data_in[3]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_3),
	.prn(vcc));
defparam \data_out_wire[3] .is_wysiwyg = "true";
defparam \data_out_wire[3] .power_up = "low";

dffeas \data_out_wire[10] (
	.clk(clock[0]),
	.d(data_in[10]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_10),
	.prn(vcc));
defparam \data_out_wire[10] .is_wysiwyg = "true";
defparam \data_out_wire[10] .power_up = "low";

dffeas \data_out_wire[2] (
	.clk(clock[0]),
	.d(data_in[2]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_2),
	.prn(vcc));
defparam \data_out_wire[2] .is_wysiwyg = "true";
defparam \data_out_wire[2] .power_up = "low";

dffeas \data_out_wire[7] (
	.clk(clock[0]),
	.d(data_in[7]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_7),
	.prn(vcc));
defparam \data_out_wire[7] .is_wysiwyg = "true";
defparam \data_out_wire[7] .power_up = "low";

dffeas \data_out_wire[6] (
	.clk(clock[0]),
	.d(data_in[6]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_6),
	.prn(vcc));
defparam \data_out_wire[6] .is_wysiwyg = "true";
defparam \data_out_wire[6] .power_up = "low";

dffeas \data_out_wire[13] (
	.clk(clock[0]),
	.d(data_in[13]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_13),
	.prn(vcc));
defparam \data_out_wire[13] .is_wysiwyg = "true";
defparam \data_out_wire[13] .power_up = "low";

dffeas \data_out_wire[14] (
	.clk(clock[0]),
	.d(data_in[14]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_14),
	.prn(vcc));
defparam \data_out_wire[14] .is_wysiwyg = "true";
defparam \data_out_wire[14] .power_up = "low";

dffeas \data_out_wire[15] (
	.clk(clock[0]),
	.d(data_in[15]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_15),
	.prn(vcc));
defparam \data_out_wire[15] .is_wysiwyg = "true";
defparam \data_out_wire[15] .power_up = "low";

dffeas \data_out_wire[12] (
	.clk(clock[0]),
	.d(data_in[12]),
	.asdata(vcc),
	.clrn(!aclr[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(data_out_wire_12),
	.prn(vcc));
defparam \data_out_wire[12] .is_wysiwyg = "true";
defparam \data_out_wire[12] .power_up = "low";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_nios2_oci (
	readdata_2,
	readdata_10,
	readdata_18,
	readdata_26,
	readdata_7,
	readdata_23,
	readdata_15,
	readdata_31,
	readdata_29,
	readdata_13,
	readdata_28,
	readdata_12,
	readdata_27,
	readdata_11,
	readdata_25,
	readdata_9,
	readdata_24,
	readdata_8,
	readdata_6,
	readdata_14,
	readdata_22,
	readdata_30,
	readdata_5,
	readdata_21,
	readdata_4,
	readdata_20,
	readdata_3,
	readdata_19,
	readdata_1,
	readdata_17,
	readdata_0,
	readdata_16,
	sr_0,
	ir_out_0,
	ir_out_1,
	d_write,
	saved_grant_0,
	waitrequest,
	mem_used_1,
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	hbreak_enabled,
	jtag_break,
	src0_valid,
	src1_valid,
	saved_grant_1,
	rf_source_valid,
	r_early_rst,
	oci_single_step_mode,
	address_nxt,
	writedata_nxt,
	debugaccess_nxt,
	byteenable_nxt,
	resetrequest,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	irf_reg_1_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	readdata_2;
output 	readdata_10;
output 	readdata_18;
output 	readdata_26;
output 	readdata_7;
output 	readdata_23;
output 	readdata_15;
output 	readdata_31;
output 	readdata_29;
output 	readdata_13;
output 	readdata_28;
output 	readdata_12;
output 	readdata_27;
output 	readdata_11;
output 	readdata_25;
output 	readdata_9;
output 	readdata_24;
output 	readdata_8;
output 	readdata_6;
output 	readdata_14;
output 	readdata_22;
output 	readdata_30;
output 	readdata_5;
output 	readdata_21;
output 	readdata_4;
output 	readdata_20;
output 	readdata_3;
output 	readdata_19;
output 	readdata_1;
output 	readdata_17;
output 	readdata_0;
output 	readdata_16;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	d_write;
input 	saved_grant_0;
output 	waitrequest;
input 	mem_used_1;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
input 	hbreak_enabled;
output 	jtag_break;
input 	src0_valid;
input 	src1_valid;
input 	saved_grant_1;
input 	rf_source_valid;
input 	r_early_rst;
output 	oci_single_step_mode;
input 	[8:0] address_nxt;
input 	[31:0] writedata_nxt;
input 	debugaccess_nxt;
input 	[3:0] byteenable_nxt;
output 	resetrequest;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[0]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[0]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[1]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[2]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[3]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[24]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[24]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[4]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[4]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[20]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[20]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[19]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[19]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[16]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[16]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[25]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[25]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[5]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[26]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[26]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[27]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[27]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[28]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[28]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[29]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[30]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[30]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[31]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[31]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[21]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[21]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[18]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[17]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[17]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[6]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[6]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[22]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[22]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[23]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[23]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[7]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[7]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[15]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[15]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[13]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[14]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[8]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[9]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[10]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[14]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[12]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[13]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[11]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_ready~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[1]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[0]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[36]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[37]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[1]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[0]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|enable_action_strobe~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[3]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[35]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_b~combout ;
wire \write~q ;
wire \read~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~1_combout ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[34]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~combout ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[25]~q ;
wire \writedata[0]~q ;
wire \address[0]~q ;
wire \address[4]~q ;
wire \address[3]~q ;
wire \address[2]~q ;
wire \address[1]~q ;
wire \address[7]~q ;
wire \address[6]~q ;
wire \address[5]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_avalon_reg|Equal0~2_combout ;
wire \debugaccess~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_avalon_reg|take_action_ocireg~0_combout ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[2]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[1]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[4]~q ;
wire \byteenable[0]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[21]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[20]~q ;
wire \write~0_combout ;
wire \write~1_combout ;
wire \write~2_combout ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[17]~q ;
wire \read~0_combout ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[3]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[2]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[5]~q ;
wire \writedata[1]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[27]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[26]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[28]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[29]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[30]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[31]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[32]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[33]~q ;
wire \writedata[3]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[19]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[18]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_error~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[6]~q ;
wire \writedata[2]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[24]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[5]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[7]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[29]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_debug|resetlatch~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[23]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[22]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[18]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[16]~q ;
wire \writedata[24]~q ;
wire \byteenable[3]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[8]~q ;
wire \writedata[4]~q ;
wire \writedata[20]~q ;
wire \byteenable[2]~q ;
wire \writedata[19]~q ;
wire \writedata[16]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ;
wire \the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_go~q ;
wire \writedata[25]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[9]~q ;
wire \writedata[5]~q ;
wire \writedata[26]~q ;
wire \writedata[27]~q ;
wire \writedata[28]~q ;
wire \writedata[29]~q ;
wire \writedata[30]~q ;
wire \writedata[31]~q ;
wire \writedata[21]~q ;
wire \writedata[18]~q ;
wire \writedata[17]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[10]~q ;
wire \writedata[10]~q ;
wire \byteenable[1]~q ;
wire \writedata[7]~q ;
wire \writedata[23]~q ;
wire \writedata[15]~q ;
wire \writedata[13]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[12]~q ;
wire \writedata[12]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[11]~q ;
wire \writedata[11]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[9]~q ;
wire \writedata[9]~q ;
wire \the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[8]~q ;
wire \writedata[8]~q ;
wire \writedata[6]~q ;
wire \writedata[14]~q ;
wire \writedata[22]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[10]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[15]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[13]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[14]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[12]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[11]~q ;
wire \readdata~0_combout ;
wire \address[8]~q ;
wire \readdata~1_combout ;
wire \readdata~2_combout ;
wire \readdata~3_combout ;


embedded_system_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper(
	.break_readreg_0(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[0]~q ),
	.MonDReg_0(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[0]~q ),
	.break_readreg_1(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[1]~q ),
	.break_readreg_2(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[2]~q ),
	.break_readreg_3(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_24(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[24]~q ),
	.MonDReg_24(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[24]~q ),
	.break_readreg_4(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[4]~q ),
	.MonDReg_4(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[4]~q ),
	.break_readreg_20(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[20]~q ),
	.MonDReg_20(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[20]~q ),
	.break_readreg_19(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[19]~q ),
	.MonDReg_19(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[19]~q ),
	.break_readreg_16(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[16]~q ),
	.MonDReg_16(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[16]~q ),
	.break_readreg_25(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[25]~q ),
	.MonDReg_25(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[25]~q ),
	.break_readreg_5(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_26(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[26]~q ),
	.MonDReg_26(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[26]~q ),
	.break_readreg_27(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[27]~q ),
	.MonDReg_27(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[27]~q ),
	.break_readreg_28(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[28]~q ),
	.MonDReg_28(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[28]~q ),
	.break_readreg_29(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[29]~q ),
	.MonDReg_30(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[30]~q ),
	.break_readreg_30(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[31]~q ),
	.MonDReg_31(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[31]~q ),
	.break_readreg_21(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[21]~q ),
	.MonDReg_21(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[21]~q ),
	.break_readreg_18(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_17(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[17]~q ),
	.MonDReg_17(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[17]~q ),
	.break_readreg_6(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[6]~q ),
	.MonDReg_6(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[6]~q ),
	.break_readreg_22(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[22]~q ),
	.MonDReg_22(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[22]~q ),
	.break_readreg_23(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[23]~q ),
	.MonDReg_23(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[23]~q ),
	.break_readreg_7(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[7]~q ),
	.MonDReg_7(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_15(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[15]~q ),
	.break_readreg_15(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[15]~q ),
	.MonDReg_13(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[14]~q ),
	.break_readreg_8(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_9(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_10(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_14(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_13(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_11(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[11]~q ),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.monitor_ready(\the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_ready~q ),
	.MonDReg_1(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[1]~q ),
	.jdo_0(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[0]~q ),
	.jdo_36(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[36]~q ),
	.jdo_37(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[37]~q ),
	.ir_1(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[1]~q ),
	.ir_0(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[3]~q ),
	.take_action_ocimem_a(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_35(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_b~combout ),
	.hbreak_enabled(hbreak_enabled),
	.take_action_ocimem_a1(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_34(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[34]~q ),
	.take_action_ocimem_a2(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~combout ),
	.jdo_25(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[25]~q ),
	.MonDReg_2(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[2]~q ),
	.jdo_1(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[1]~q ),
	.jdo_4(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[4]~q ),
	.jdo_21(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[20]~q ),
	.jdo_17(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[17]~q ),
	.MonDReg_3(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[3]~q ),
	.jdo_2(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[2]~q ),
	.jdo_5(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[5]~q ),
	.jdo_27(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[27]~q ),
	.jdo_26(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[26]~q ),
	.jdo_28(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[28]~q ),
	.jdo_29(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[29]~q ),
	.jdo_30(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[30]~q ),
	.jdo_31(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[31]~q ),
	.jdo_32(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[32]~q ),
	.jdo_33(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[33]~q ),
	.jdo_19(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[18]~q ),
	.monitor_error(\the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_error~q ),
	.jdo_6(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[6]~q ),
	.jdo_24(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[24]~q ),
	.MonDReg_5(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[5]~q ),
	.jdo_7(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[7]~q ),
	.MonDReg_29(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[29]~q ),
	.resetlatch(\the_embedded_system_nios2_qsys_0_nios2_oci_debug|resetlatch~q ),
	.jdo_23(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[22]~q ),
	.MonDReg_18(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[18]~q ),
	.jdo_16(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[16]~q ),
	.jdo_8(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[8]~q ),
	.jdo_9(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[9]~q ),
	.MonDReg_10(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[10]~q ),
	.MonDReg_12(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[12]~q ),
	.MonDReg_11(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[11]~q ),
	.MonDReg_9(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[9]~q ),
	.MonDReg_8(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[8]~q ),
	.jdo_10(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[10]~q ),
	.jdo_15(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[15]~q ),
	.jdo_13(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[13]~q ),
	.jdo_14(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[14]~q ),
	.jdo_12(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[12]~q ),
	.jdo_11(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[11]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_nios2_oci_break the_embedded_system_nios2_qsys_0_nios2_oci_break(
	.break_readreg_0(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[0]~q ),
	.break_readreg_1(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[1]~q ),
	.break_readreg_2(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[2]~q ),
	.break_readreg_3(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[3]~q ),
	.break_readreg_24(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[24]~q ),
	.break_readreg_4(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[4]~q ),
	.break_readreg_20(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[20]~q ),
	.break_readreg_19(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[19]~q ),
	.break_readreg_16(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[16]~q ),
	.break_readreg_25(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[25]~q ),
	.break_readreg_5(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[5]~q ),
	.break_readreg_26(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[26]~q ),
	.break_readreg_27(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[27]~q ),
	.break_readreg_28(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[28]~q ),
	.break_readreg_29(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[29]~q ),
	.break_readreg_30(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[30]~q ),
	.break_readreg_31(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[31]~q ),
	.break_readreg_21(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[21]~q ),
	.break_readreg_18(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[18]~q ),
	.break_readreg_17(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[17]~q ),
	.break_readreg_6(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[6]~q ),
	.break_readreg_22(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[22]~q ),
	.break_readreg_23(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[23]~q ),
	.break_readreg_7(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[7]~q ),
	.break_readreg_15(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[15]~q ),
	.break_readreg_8(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[8]~q ),
	.break_readreg_9(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[9]~q ),
	.break_readreg_10(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[10]~q ),
	.break_readreg_14(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[14]~q ),
	.break_readreg_12(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[12]~q ),
	.break_readreg_13(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[13]~q ),
	.break_readreg_11(\the_embedded_system_nios2_qsys_0_nios2_oci_break|break_readreg[11]~q ),
	.jdo_0(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[0]~q ),
	.jdo_36(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[36]~q ),
	.jdo_37(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[37]~q ),
	.ir_1(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[1]~q ),
	.ir_0(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|ir[0]~q ),
	.enable_action_strobe(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|enable_action_strobe~q ),
	.jdo_3(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[3]~q ),
	.jdo_25(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[25]~q ),
	.jdo_1(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[1]~q ),
	.jdo_4(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[4]~q ),
	.jdo_21(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[20]~q ),
	.jdo_17(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[17]~q ),
	.jdo_2(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[2]~q ),
	.jdo_5(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[5]~q ),
	.jdo_27(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[27]~q ),
	.jdo_26(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[26]~q ),
	.jdo_28(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[28]~q ),
	.jdo_29(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[29]~q ),
	.jdo_30(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[30]~q ),
	.jdo_31(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[31]~q ),
	.jdo_19(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[18]~q ),
	.jdo_6(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[6]~q ),
	.jdo_24(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[24]~q ),
	.jdo_7(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[7]~q ),
	.jdo_23(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[22]~q ),
	.jdo_16(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[16]~q ),
	.jdo_8(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[8]~q ),
	.jdo_9(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[9]~q ),
	.jdo_10(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[10]~q ),
	.jdo_15(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[15]~q ),
	.jdo_13(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[13]~q ),
	.jdo_14(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[14]~q ),
	.jdo_12(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[12]~q ),
	.jdo_11(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[11]~q ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_nios2_avalon_reg the_embedded_system_nios2_qsys_0_nios2_avalon_reg(
	.hq3myc14108phmpo7y7qmhbp98hy0vq(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.address_0(\address[0]~q ),
	.address_4(\address[4]~q ),
	.address_3(\address[3]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.Equal0(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|Equal0~2_combout ),
	.debugaccess(\debugaccess~q ),
	.take_action_ocireg(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.oci_single_step_mode1(oci_single_step_mode),
	.writedata_3(\writedata[3]~q ),
	.oci_reg_readdata(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_nios2_ocimem the_embedded_system_nios2_qsys_0_nios2_ocimem(
	.MonDReg_0(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[0]~q ),
	.q_a_0(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.q_a_1(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.q_a_2(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.MonDReg_24(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[24]~q ),
	.MonDReg_4(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[4]~q ),
	.q_a_3(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.MonDReg_20(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[20]~q ),
	.MonDReg_19(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[19]~q ),
	.MonDReg_16(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[16]~q ),
	.MonDReg_25(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[25]~q ),
	.q_a_24(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.q_a_4(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.MonDReg_26(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[26]~q ),
	.MonDReg_27(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[27]~q ),
	.MonDReg_28(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[28]~q ),
	.MonDReg_30(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[30]~q ),
	.MonDReg_31(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[31]~q ),
	.MonDReg_21(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[21]~q ),
	.q_a_20(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.q_a_19(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.MonDReg_17(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[17]~q ),
	.q_a_16(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.q_a_25(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.MonDReg_6(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[6]~q ),
	.q_a_5(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.q_a_26(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.q_a_27(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.q_a_28(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.q_a_29(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.q_a_30(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.q_a_31(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.MonDReg_22(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[22]~q ),
	.q_a_21(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.q_a_18(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.q_a_17(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.q_a_10(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.q_a_7(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.q_a_23(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.q_a_15(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.q_a_13(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.q_a_12(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.q_a_11(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.q_a_9(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.q_a_8(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.q_a_6(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.q_a_14(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.q_a_22(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.MonDReg_23(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[23]~q ),
	.MonDReg_7(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[7]~q ),
	.MonDReg_15(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[15]~q ),
	.MonDReg_13(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[13]~q ),
	.MonDReg_14(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[14]~q ),
	.waitrequest1(waitrequest),
	.MonDReg_1(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[1]~q ),
	.jdo_3(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[3]~q ),
	.take_action_ocimem_a(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~0_combout ),
	.jdo_35(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[35]~q ),
	.take_action_ocimem_b(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_b~combout ),
	.write(\write~q ),
	.address_8(\address[8]~q ),
	.read(\read~q ),
	.take_action_ocimem_a1(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_34(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[34]~q ),
	.take_action_ocimem_a2(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~combout ),
	.jdo_25(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.address_0(\address[0]~q ),
	.address_4(\address[4]~q ),
	.address_3(\address[3]~q ),
	.address_2(\address[2]~q ),
	.address_1(\address[1]~q ),
	.address_7(\address[7]~q ),
	.address_6(\address[6]~q ),
	.address_5(\address[5]~q ),
	.debugaccess(\debugaccess~q ),
	.MonDReg_2(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[2]~q ),
	.jdo_4(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[4]~q ),
	.r_early_rst(r_early_rst),
	.byteenable_0(\byteenable[0]~q ),
	.jdo_21(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[20]~q ),
	.jdo_17(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[17]~q ),
	.MonDReg_3(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[3]~q ),
	.jdo_5(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[5]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_27(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[27]~q ),
	.jdo_26(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[26]~q ),
	.jdo_28(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[28]~q ),
	.jdo_29(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[29]~q ),
	.jdo_30(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[30]~q ),
	.jdo_31(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[31]~q ),
	.jdo_32(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[32]~q ),
	.jdo_33(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[33]~q ),
	.writedata_3(\writedata[3]~q ),
	.jdo_19(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[18]~q ),
	.jdo_6(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[6]~q ),
	.writedata_2(\writedata[2]~q ),
	.jdo_24(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[24]~q ),
	.MonDReg_5(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[5]~q ),
	.jdo_7(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[7]~q ),
	.MonDReg_29(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[29]~q ),
	.jdo_23(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[22]~q ),
	.MonDReg_18(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[18]~q ),
	.jdo_16(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[16]~q ),
	.writedata_24(\writedata[24]~q ),
	.byteenable_3(\byteenable[3]~q ),
	.jdo_8(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[8]~q ),
	.writedata_4(\writedata[4]~q ),
	.writedata_20(\writedata[20]~q ),
	.byteenable_2(\byteenable[2]~q ),
	.writedata_19(\writedata[19]~q ),
	.writedata_16(\writedata[16]~q ),
	.writedata_25(\writedata[25]~q ),
	.jdo_9(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[9]~q ),
	.writedata_5(\writedata[5]~q ),
	.writedata_26(\writedata[26]~q ),
	.writedata_27(\writedata[27]~q ),
	.writedata_28(\writedata[28]~q ),
	.writedata_29(\writedata[29]~q ),
	.writedata_30(\writedata[30]~q ),
	.writedata_31(\writedata[31]~q ),
	.writedata_21(\writedata[21]~q ),
	.writedata_18(\writedata[18]~q ),
	.writedata_17(\writedata[17]~q ),
	.MonDReg_10(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[10]~q ),
	.writedata_10(\writedata[10]~q ),
	.byteenable_1(\byteenable[1]~q ),
	.writedata_7(\writedata[7]~q ),
	.writedata_23(\writedata[23]~q ),
	.writedata_15(\writedata[15]~q ),
	.writedata_13(\writedata[13]~q ),
	.MonDReg_12(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[12]~q ),
	.writedata_12(\writedata[12]~q ),
	.MonDReg_11(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[11]~q ),
	.writedata_11(\writedata[11]~q ),
	.MonDReg_9(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[9]~q ),
	.writedata_9(\writedata[9]~q ),
	.MonDReg_8(\the_embedded_system_nios2_qsys_0_nios2_ocimem|MonDReg[8]~q ),
	.writedata_8(\writedata[8]~q ),
	.writedata_6(\writedata[6]~q ),
	.writedata_14(\writedata[14]~q ),
	.writedata_22(\writedata[22]~q ),
	.jdo_10(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[10]~q ),
	.jdo_15(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[15]~q ),
	.jdo_13(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[13]~q ),
	.jdo_14(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[14]~q ),
	.jdo_12(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[12]~q ),
	.jdo_11(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[11]~q ),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_nios2_oci_debug the_embedded_system_nios2_qsys_0_nios2_oci_debug(
	.hq3myc14108phmpo7y7qmhbp98hy0vq(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.monitor_ready1(\the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_ready~q ),
	.jtag_break1(jtag_break),
	.take_action_ocimem_a(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~1_combout ),
	.jdo_34(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[34]~q ),
	.take_action_ocimem_a1(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|take_action_ocimem_a~combout ),
	.jdo_25(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[25]~q ),
	.writedata_0(\writedata[0]~q ),
	.take_action_ocireg(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|take_action_ocireg~0_combout ),
	.jdo_21(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[21]~q ),
	.jdo_20(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[20]~q ),
	.writedata_1(\writedata[1]~q ),
	.jdo_19(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[19]~q ),
	.jdo_18(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[18]~q ),
	.monitor_error1(\the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_error~q ),
	.resetrequest1(resetrequest),
	.jdo_24(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[24]~q ),
	.resetlatch1(\the_embedded_system_nios2_qsys_0_nios2_oci_debug|resetlatch~q ),
	.jdo_23(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[23]~q ),
	.jdo_22(\the_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper|the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk|jdo[22]~q ),
	.monitor_go1(\the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_go~q ),
	.state_1(state_1),
	.clk_clk(clk_clk));

dffeas write(
	.clk(clk_clk),
	.d(\write~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\write~q ),
	.prn(vcc));
defparam write.is_wysiwyg = "true";
defparam write.power_up = "low";

dffeas read(
	.clk(clk_clk),
	.d(\read~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\read~q ),
	.prn(vcc));
defparam read.is_wysiwyg = "true";
defparam read.power_up = "low";

dffeas \writedata[0] (
	.clk(clk_clk),
	.d(writedata_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[0]~q ),
	.prn(vcc));
defparam \writedata[0] .is_wysiwyg = "true";
defparam \writedata[0] .power_up = "low";

dffeas \address[0] (
	.clk(clk_clk),
	.d(address_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[0]~q ),
	.prn(vcc));
defparam \address[0] .is_wysiwyg = "true";
defparam \address[0] .power_up = "low";

dffeas \address[4] (
	.clk(clk_clk),
	.d(address_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[4]~q ),
	.prn(vcc));
defparam \address[4] .is_wysiwyg = "true";
defparam \address[4] .power_up = "low";

dffeas \address[3] (
	.clk(clk_clk),
	.d(address_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[3]~q ),
	.prn(vcc));
defparam \address[3] .is_wysiwyg = "true";
defparam \address[3] .power_up = "low";

dffeas \address[2] (
	.clk(clk_clk),
	.d(address_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[2]~q ),
	.prn(vcc));
defparam \address[2] .is_wysiwyg = "true";
defparam \address[2] .power_up = "low";

dffeas \address[1] (
	.clk(clk_clk),
	.d(address_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[1]~q ),
	.prn(vcc));
defparam \address[1] .is_wysiwyg = "true";
defparam \address[1] .power_up = "low";

dffeas \address[7] (
	.clk(clk_clk),
	.d(address_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[7]~q ),
	.prn(vcc));
defparam \address[7] .is_wysiwyg = "true";
defparam \address[7] .power_up = "low";

dffeas \address[6] (
	.clk(clk_clk),
	.d(address_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[6]~q ),
	.prn(vcc));
defparam \address[6] .is_wysiwyg = "true";
defparam \address[6] .power_up = "low";

dffeas \address[5] (
	.clk(clk_clk),
	.d(address_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[5]~q ),
	.prn(vcc));
defparam \address[5] .is_wysiwyg = "true";
defparam \address[5] .power_up = "low";

dffeas debugaccess(
	.clk(clk_clk),
	.d(debugaccess_nxt),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\debugaccess~q ),
	.prn(vcc));
defparam debugaccess.is_wysiwyg = "true";
defparam debugaccess.power_up = "low";

dffeas \byteenable[0] (
	.clk(clk_clk),
	.d(byteenable_nxt[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[0]~q ),
	.prn(vcc));
defparam \byteenable[0] .is_wysiwyg = "true";
defparam \byteenable[0] .power_up = "low";

cyclonev_lcell_comb \write~0 (
	.dataa(!d_write),
	.datab(!mem_used_1),
	.datac(!\write~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~0 .extended_lut = "off";
defparam \write~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \write~0 .shared_arith = "off";

cyclonev_lcell_comb \write~1 (
	.dataa(!saved_grant_0),
	.datab(!src0_valid),
	.datac(!src1_valid),
	.datad(!saved_grant_1),
	.datae(!\write~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~1 .extended_lut = "off";
defparam \write~1 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \write~1 .shared_arith = "off";

cyclonev_lcell_comb \write~2 (
	.dataa(!waitrequest),
	.datab(!\write~q ),
	.datac(!\write~1_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\write~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \write~2 .extended_lut = "off";
defparam \write~2 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \write~2 .shared_arith = "off";

cyclonev_lcell_comb \read~0 (
	.dataa(!waitrequest),
	.datab(!mem_used_1),
	.datac(!\read~q ),
	.datad(!rf_source_valid),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\read~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \read~0 .extended_lut = "off";
defparam \read~0 .lut_mask = 64'hC5FFC5FFC5FFC5FF;
defparam \read~0 .shared_arith = "off";

dffeas \writedata[1] (
	.clk(clk_clk),
	.d(writedata_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[1]~q ),
	.prn(vcc));
defparam \writedata[1] .is_wysiwyg = "true";
defparam \writedata[1] .power_up = "low";

dffeas \writedata[3] (
	.clk(clk_clk),
	.d(writedata_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[3]~q ),
	.prn(vcc));
defparam \writedata[3] .is_wysiwyg = "true";
defparam \writedata[3] .power_up = "low";

dffeas \writedata[2] (
	.clk(clk_clk),
	.d(writedata_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[2]~q ),
	.prn(vcc));
defparam \writedata[2] .is_wysiwyg = "true";
defparam \writedata[2] .power_up = "low";

dffeas \writedata[24] (
	.clk(clk_clk),
	.d(writedata_nxt[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[24]~q ),
	.prn(vcc));
defparam \writedata[24] .is_wysiwyg = "true";
defparam \writedata[24] .power_up = "low";

dffeas \byteenable[3] (
	.clk(clk_clk),
	.d(byteenable_nxt[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[3]~q ),
	.prn(vcc));
defparam \byteenable[3] .is_wysiwyg = "true";
defparam \byteenable[3] .power_up = "low";

dffeas \writedata[4] (
	.clk(clk_clk),
	.d(writedata_nxt[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[4]~q ),
	.prn(vcc));
defparam \writedata[4] .is_wysiwyg = "true";
defparam \writedata[4] .power_up = "low";

dffeas \writedata[20] (
	.clk(clk_clk),
	.d(writedata_nxt[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[20]~q ),
	.prn(vcc));
defparam \writedata[20] .is_wysiwyg = "true";
defparam \writedata[20] .power_up = "low";

dffeas \byteenable[2] (
	.clk(clk_clk),
	.d(byteenable_nxt[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[2]~q ),
	.prn(vcc));
defparam \byteenable[2] .is_wysiwyg = "true";
defparam \byteenable[2] .power_up = "low";

dffeas \writedata[19] (
	.clk(clk_clk),
	.d(writedata_nxt[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[19]~q ),
	.prn(vcc));
defparam \writedata[19] .is_wysiwyg = "true";
defparam \writedata[19] .power_up = "low";

dffeas \writedata[16] (
	.clk(clk_clk),
	.d(writedata_nxt[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[16]~q ),
	.prn(vcc));
defparam \writedata[16] .is_wysiwyg = "true";
defparam \writedata[16] .power_up = "low";

dffeas \writedata[25] (
	.clk(clk_clk),
	.d(writedata_nxt[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[25]~q ),
	.prn(vcc));
defparam \writedata[25] .is_wysiwyg = "true";
defparam \writedata[25] .power_up = "low";

dffeas \writedata[5] (
	.clk(clk_clk),
	.d(writedata_nxt[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[5]~q ),
	.prn(vcc));
defparam \writedata[5] .is_wysiwyg = "true";
defparam \writedata[5] .power_up = "low";

dffeas \writedata[26] (
	.clk(clk_clk),
	.d(writedata_nxt[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[26]~q ),
	.prn(vcc));
defparam \writedata[26] .is_wysiwyg = "true";
defparam \writedata[26] .power_up = "low";

dffeas \writedata[27] (
	.clk(clk_clk),
	.d(writedata_nxt[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[27]~q ),
	.prn(vcc));
defparam \writedata[27] .is_wysiwyg = "true";
defparam \writedata[27] .power_up = "low";

dffeas \writedata[28] (
	.clk(clk_clk),
	.d(writedata_nxt[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[28]~q ),
	.prn(vcc));
defparam \writedata[28] .is_wysiwyg = "true";
defparam \writedata[28] .power_up = "low";

dffeas \writedata[29] (
	.clk(clk_clk),
	.d(writedata_nxt[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[29]~q ),
	.prn(vcc));
defparam \writedata[29] .is_wysiwyg = "true";
defparam \writedata[29] .power_up = "low";

dffeas \writedata[30] (
	.clk(clk_clk),
	.d(writedata_nxt[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[30]~q ),
	.prn(vcc));
defparam \writedata[30] .is_wysiwyg = "true";
defparam \writedata[30] .power_up = "low";

dffeas \writedata[31] (
	.clk(clk_clk),
	.d(writedata_nxt[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[31]~q ),
	.prn(vcc));
defparam \writedata[31] .is_wysiwyg = "true";
defparam \writedata[31] .power_up = "low";

dffeas \writedata[21] (
	.clk(clk_clk),
	.d(writedata_nxt[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[21]~q ),
	.prn(vcc));
defparam \writedata[21] .is_wysiwyg = "true";
defparam \writedata[21] .power_up = "low";

dffeas \writedata[18] (
	.clk(clk_clk),
	.d(writedata_nxt[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[18]~q ),
	.prn(vcc));
defparam \writedata[18] .is_wysiwyg = "true";
defparam \writedata[18] .power_up = "low";

dffeas \writedata[17] (
	.clk(clk_clk),
	.d(writedata_nxt[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[17]~q ),
	.prn(vcc));
defparam \writedata[17] .is_wysiwyg = "true";
defparam \writedata[17] .power_up = "low";

dffeas \writedata[10] (
	.clk(clk_clk),
	.d(writedata_nxt[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[10]~q ),
	.prn(vcc));
defparam \writedata[10] .is_wysiwyg = "true";
defparam \writedata[10] .power_up = "low";

dffeas \byteenable[1] (
	.clk(clk_clk),
	.d(byteenable_nxt[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\byteenable[1]~q ),
	.prn(vcc));
defparam \byteenable[1] .is_wysiwyg = "true";
defparam \byteenable[1] .power_up = "low";

dffeas \writedata[7] (
	.clk(clk_clk),
	.d(writedata_nxt[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[7]~q ),
	.prn(vcc));
defparam \writedata[7] .is_wysiwyg = "true";
defparam \writedata[7] .power_up = "low";

dffeas \writedata[23] (
	.clk(clk_clk),
	.d(writedata_nxt[23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[23]~q ),
	.prn(vcc));
defparam \writedata[23] .is_wysiwyg = "true";
defparam \writedata[23] .power_up = "low";

dffeas \writedata[15] (
	.clk(clk_clk),
	.d(writedata_nxt[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[15]~q ),
	.prn(vcc));
defparam \writedata[15] .is_wysiwyg = "true";
defparam \writedata[15] .power_up = "low";

dffeas \writedata[13] (
	.clk(clk_clk),
	.d(writedata_nxt[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[13]~q ),
	.prn(vcc));
defparam \writedata[13] .is_wysiwyg = "true";
defparam \writedata[13] .power_up = "low";

dffeas \writedata[12] (
	.clk(clk_clk),
	.d(writedata_nxt[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[12]~q ),
	.prn(vcc));
defparam \writedata[12] .is_wysiwyg = "true";
defparam \writedata[12] .power_up = "low";

dffeas \writedata[11] (
	.clk(clk_clk),
	.d(writedata_nxt[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[11]~q ),
	.prn(vcc));
defparam \writedata[11] .is_wysiwyg = "true";
defparam \writedata[11] .power_up = "low";

dffeas \writedata[9] (
	.clk(clk_clk),
	.d(writedata_nxt[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[9]~q ),
	.prn(vcc));
defparam \writedata[9] .is_wysiwyg = "true";
defparam \writedata[9] .power_up = "low";

dffeas \writedata[8] (
	.clk(clk_clk),
	.d(writedata_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[8]~q ),
	.prn(vcc));
defparam \writedata[8] .is_wysiwyg = "true";
defparam \writedata[8] .power_up = "low";

dffeas \writedata[6] (
	.clk(clk_clk),
	.d(writedata_nxt[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[6]~q ),
	.prn(vcc));
defparam \writedata[6] .is_wysiwyg = "true";
defparam \writedata[6] .power_up = "low";

dffeas \writedata[14] (
	.clk(clk_clk),
	.d(writedata_nxt[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[14]~q ),
	.prn(vcc));
defparam \writedata[14] .is_wysiwyg = "true";
defparam \writedata[14] .power_up = "low";

dffeas \writedata[22] (
	.clk(clk_clk),
	.d(writedata_nxt[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\writedata[22]~q ),
	.prn(vcc));
defparam \writedata[22] .is_wysiwyg = "true";
defparam \writedata[22] .power_up = "low";

dffeas \readdata[2] (
	.clk(clk_clk),
	.d(\readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[2] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_2),
	.prn(vcc));
defparam \readdata[2] .is_wysiwyg = "true";
defparam \readdata[2] .power_up = "low";

dffeas \readdata[10] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[10] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_10),
	.prn(vcc));
defparam \readdata[10] .is_wysiwyg = "true";
defparam \readdata[10] .power_up = "low";

dffeas \readdata[18] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[18] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_18),
	.prn(vcc));
defparam \readdata[18] .is_wysiwyg = "true";
defparam \readdata[18] .power_up = "low";

dffeas \readdata[26] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[26] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_26),
	.prn(vcc));
defparam \readdata[26] .is_wysiwyg = "true";
defparam \readdata[26] .power_up = "low";

dffeas \readdata[7] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[7] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_7),
	.prn(vcc));
defparam \readdata[7] .is_wysiwyg = "true";
defparam \readdata[7] .power_up = "low";

dffeas \readdata[23] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[23] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_23),
	.prn(vcc));
defparam \readdata[23] .is_wysiwyg = "true";
defparam \readdata[23] .power_up = "low";

dffeas \readdata[15] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[15] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_15),
	.prn(vcc));
defparam \readdata[15] .is_wysiwyg = "true";
defparam \readdata[15] .power_up = "low";

dffeas \readdata[31] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[31] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_31),
	.prn(vcc));
defparam \readdata[31] .is_wysiwyg = "true";
defparam \readdata[31] .power_up = "low";

dffeas \readdata[29] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[29] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_29),
	.prn(vcc));
defparam \readdata[29] .is_wysiwyg = "true";
defparam \readdata[29] .power_up = "low";

dffeas \readdata[13] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[13] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_13),
	.prn(vcc));
defparam \readdata[13] .is_wysiwyg = "true";
defparam \readdata[13] .power_up = "low";

dffeas \readdata[28] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[28] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_28),
	.prn(vcc));
defparam \readdata[28] .is_wysiwyg = "true";
defparam \readdata[28] .power_up = "low";

dffeas \readdata[12] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[12] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_12),
	.prn(vcc));
defparam \readdata[12] .is_wysiwyg = "true";
defparam \readdata[12] .power_up = "low";

dffeas \readdata[27] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[27] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_27),
	.prn(vcc));
defparam \readdata[27] .is_wysiwyg = "true";
defparam \readdata[27] .power_up = "low";

dffeas \readdata[11] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[11] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_11),
	.prn(vcc));
defparam \readdata[11] .is_wysiwyg = "true";
defparam \readdata[11] .power_up = "low";

dffeas \readdata[25] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[25] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_25),
	.prn(vcc));
defparam \readdata[25] .is_wysiwyg = "true";
defparam \readdata[25] .power_up = "low";

dffeas \readdata[9] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[9] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_9),
	.prn(vcc));
defparam \readdata[9] .is_wysiwyg = "true";
defparam \readdata[9] .power_up = "low";

dffeas \readdata[24] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[24] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_24),
	.prn(vcc));
defparam \readdata[24] .is_wysiwyg = "true";
defparam \readdata[24] .power_up = "low";

dffeas \readdata[8] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[8] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_8),
	.prn(vcc));
defparam \readdata[8] .is_wysiwyg = "true";
defparam \readdata[8] .power_up = "low";

dffeas \readdata[6] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[6] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_6),
	.prn(vcc));
defparam \readdata[6] .is_wysiwyg = "true";
defparam \readdata[6] .power_up = "low";

dffeas \readdata[14] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[14] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_14),
	.prn(vcc));
defparam \readdata[14] .is_wysiwyg = "true";
defparam \readdata[14] .power_up = "low";

dffeas \readdata[22] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[22] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_22),
	.prn(vcc));
defparam \readdata[22] .is_wysiwyg = "true";
defparam \readdata[22] .power_up = "low";

dffeas \readdata[30] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[30] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_30),
	.prn(vcc));
defparam \readdata[30] .is_wysiwyg = "true";
defparam \readdata[30] .power_up = "low";

dffeas \readdata[5] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[5] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_5),
	.prn(vcc));
defparam \readdata[5] .is_wysiwyg = "true";
defparam \readdata[5] .power_up = "low";

dffeas \readdata[21] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[21] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_21),
	.prn(vcc));
defparam \readdata[21] .is_wysiwyg = "true";
defparam \readdata[21] .power_up = "low";

dffeas \readdata[4] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[4] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_4),
	.prn(vcc));
defparam \readdata[4] .is_wysiwyg = "true";
defparam \readdata[4] .power_up = "low";

dffeas \readdata[20] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[20] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_20),
	.prn(vcc));
defparam \readdata[20] .is_wysiwyg = "true";
defparam \readdata[20] .power_up = "low";

dffeas \readdata[3] (
	.clk(clk_clk),
	.d(\readdata~1_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[3] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_3),
	.prn(vcc));
defparam \readdata[3] .is_wysiwyg = "true";
defparam \readdata[3] .power_up = "low";

dffeas \readdata[19] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[19] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_19),
	.prn(vcc));
defparam \readdata[19] .is_wysiwyg = "true";
defparam \readdata[19] .power_up = "low";

dffeas \readdata[1] (
	.clk(clk_clk),
	.d(\readdata~2_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[1] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_1),
	.prn(vcc));
defparam \readdata[1] .is_wysiwyg = "true";
defparam \readdata[1] .power_up = "low";

dffeas \readdata[17] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[17] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_17),
	.prn(vcc));
defparam \readdata[17] .is_wysiwyg = "true";
defparam \readdata[17] .power_up = "low";

dffeas \readdata[0] (
	.clk(clk_clk),
	.d(\readdata~3_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[0] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_0),
	.prn(vcc));
defparam \readdata[0] .is_wysiwyg = "true";
defparam \readdata[0] .power_up = "low";

dffeas \readdata[16] (
	.clk(clk_clk),
	.d(\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.asdata(\the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram|the_altsyncram|auto_generated|q_a[16] ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\address[8]~q ),
	.ena(vcc),
	.q(readdata_16),
	.prn(vcc));
defparam \readdata[16] .is_wysiwyg = "true";
defparam \readdata[16] .power_up = "low";

cyclonev_lcell_comb \readdata~0 (
	.dataa(!\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|Equal0~2_combout ),
	.datab(!\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.datac(!\the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_go~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~0 .extended_lut = "off";
defparam \readdata~0 .lut_mask = 64'h2727272727272727;
defparam \readdata~0 .shared_arith = "off";

dffeas \address[8] (
	.clk(clk_clk),
	.d(address_nxt[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\address[8]~q ),
	.prn(vcc));
defparam \address[8] .is_wysiwyg = "true";
defparam \address[8] .power_up = "low";

cyclonev_lcell_comb \readdata~1 (
	.dataa(!\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|Equal0~2_combout ),
	.datab(!oci_single_step_mode),
	.datac(!\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~1 .extended_lut = "off";
defparam \readdata~1 .lut_mask = 64'h2727272727272727;
defparam \readdata~1 .shared_arith = "off";

cyclonev_lcell_comb \readdata~2 (
	.dataa(!\the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_ready~q ),
	.datab(!\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|Equal0~2_combout ),
	.datac(!\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~2 .extended_lut = "off";
defparam \readdata~2 .lut_mask = 64'h4747474747474747;
defparam \readdata~2 .shared_arith = "off";

cyclonev_lcell_comb \readdata~3 (
	.dataa(!\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|Equal0~2_combout ),
	.datab(!\the_embedded_system_nios2_qsys_0_nios2_oci_debug|monitor_error~q ),
	.datac(!\the_embedded_system_nios2_qsys_0_nios2_avalon_reg|oci_reg_readdata~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\readdata~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \readdata~3 .extended_lut = "off";
defparam \readdata~3 .lut_mask = 64'h2727272727272727;
defparam \readdata~3 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_jtag_debug_module_wrapper (
	break_readreg_0,
	MonDReg_0,
	break_readreg_1,
	break_readreg_2,
	break_readreg_3,
	break_readreg_24,
	MonDReg_24,
	break_readreg_4,
	MonDReg_4,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	break_readreg_16,
	MonDReg_16,
	break_readreg_25,
	MonDReg_25,
	break_readreg_5,
	break_readreg_26,
	MonDReg_26,
	break_readreg_27,
	MonDReg_27,
	break_readreg_28,
	MonDReg_28,
	break_readreg_29,
	MonDReg_30,
	break_readreg_30,
	break_readreg_31,
	MonDReg_31,
	break_readreg_21,
	MonDReg_21,
	break_readreg_18,
	break_readreg_17,
	MonDReg_17,
	break_readreg_6,
	MonDReg_6,
	break_readreg_22,
	MonDReg_22,
	break_readreg_23,
	MonDReg_23,
	break_readreg_7,
	MonDReg_7,
	MonDReg_15,
	break_readreg_15,
	MonDReg_13,
	MonDReg_14,
	break_readreg_8,
	break_readreg_9,
	break_readreg_10,
	break_readreg_14,
	break_readreg_12,
	break_readreg_13,
	break_readreg_11,
	sr_0,
	ir_out_0,
	ir_out_1,
	monitor_ready,
	MonDReg_1,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe,
	jdo_3,
	take_action_ocimem_a,
	jdo_35,
	take_action_ocimem_b,
	hbreak_enabled,
	take_action_ocimem_a1,
	jdo_34,
	take_action_ocimem_a2,
	jdo_25,
	MonDReg_2,
	jdo_1,
	jdo_4,
	jdo_21,
	jdo_20,
	jdo_17,
	MonDReg_3,
	jdo_2,
	jdo_5,
	jdo_27,
	jdo_26,
	jdo_28,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_19,
	jdo_18,
	monitor_error,
	jdo_6,
	jdo_24,
	MonDReg_5,
	jdo_7,
	MonDReg_29,
	resetlatch,
	jdo_23,
	jdo_22,
	MonDReg_18,
	jdo_16,
	jdo_8,
	jdo_9,
	MonDReg_10,
	MonDReg_12,
	MonDReg_11,
	MonDReg_9,
	MonDReg_8,
	jdo_10,
	jdo_15,
	jdo_13,
	jdo_14,
	jdo_12,
	jdo_11,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	irf_reg_0_1,
	irf_reg_1_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	break_readreg_0;
input 	MonDReg_0;
input 	break_readreg_1;
input 	break_readreg_2;
input 	break_readreg_3;
input 	break_readreg_24;
input 	MonDReg_24;
input 	break_readreg_4;
input 	MonDReg_4;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_5;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_29;
input 	MonDReg_30;
input 	break_readreg_30;
input 	break_readreg_31;
input 	MonDReg_31;
input 	break_readreg_21;
input 	MonDReg_21;
input 	break_readreg_18;
input 	break_readreg_17;
input 	MonDReg_17;
input 	break_readreg_6;
input 	MonDReg_6;
input 	break_readreg_22;
input 	MonDReg_22;
input 	break_readreg_23;
input 	MonDReg_23;
input 	break_readreg_7;
input 	MonDReg_7;
input 	MonDReg_15;
input 	break_readreg_15;
input 	MonDReg_13;
input 	MonDReg_14;
input 	break_readreg_8;
input 	break_readreg_9;
input 	break_readreg_10;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_13;
input 	break_readreg_11;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	monitor_ready;
input 	MonDReg_1;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe;
output 	jdo_3;
output 	take_action_ocimem_a;
output 	jdo_35;
output 	take_action_ocimem_b;
input 	hbreak_enabled;
output 	take_action_ocimem_a1;
output 	jdo_34;
output 	take_action_ocimem_a2;
output 	jdo_25;
input 	MonDReg_2;
output 	jdo_1;
output 	jdo_4;
output 	jdo_21;
output 	jdo_20;
output 	jdo_17;
input 	MonDReg_3;
output 	jdo_2;
output 	jdo_5;
output 	jdo_27;
output 	jdo_26;
output 	jdo_28;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
output 	jdo_19;
output 	jdo_18;
input 	monitor_error;
output 	jdo_6;
output 	jdo_24;
input 	MonDReg_5;
output 	jdo_7;
input 	MonDReg_29;
input 	resetlatch;
output 	jdo_23;
output 	jdo_22;
input 	MonDReg_18;
output 	jdo_16;
output 	jdo_8;
output 	jdo_9;
input 	MonDReg_10;
input 	MonDReg_12;
input 	MonDReg_11;
input 	MonDReg_9;
input 	MonDReg_8;
output 	jdo_10;
output 	jdo_15;
output 	jdo_13;
output 	jdo_14;
output 	jdo_12;
output 	jdo_11;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[1]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[2]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[3]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[4]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[25]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[5]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[21]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[20]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[17]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[26]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[6]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[27]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[28]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[29]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[30]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[32]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[22]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[19]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[18]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[23]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[24]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[8]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[16]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[9]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[10]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[11]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[13]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[14]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[12]~q ;
wire \embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_sdr~0_combout ;
wire \embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_uir~combout ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[36]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[37]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[35]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[34]~q ;
wire \embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_cdr~combout ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[31]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[33]~q ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[7]~q ;
wire \embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_udr~0_combout ;
wire \the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[15]~q ;


embedded_system_sld_virtual_jtag_basic_1 embedded_system_nios2_qsys_0_jtag_debug_module_phy(
	.virtual_state_sdr(\embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir1(\embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_uir~combout ),
	.virtual_state_cdr1(\embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_cdr~combout ),
	.virtual_state_udr(\embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_udr~0_combout ),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8));

embedded_system_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk the_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk(
	.sr_1(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[1]~q ),
	.sr_2(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[2]~q ),
	.sr_3(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[3]~q ),
	.sr_4(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[4]~q ),
	.sr_25(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[25]~q ),
	.sr_5(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[5]~q ),
	.sr_21(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[21]~q ),
	.sr_20(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[20]~q ),
	.sr_17(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[17]~q ),
	.sr_26(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[26]~q ),
	.sr_6(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[6]~q ),
	.sr_27(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[27]~q ),
	.sr_28(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[28]~q ),
	.sr_29(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[29]~q ),
	.sr_30(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[30]~q ),
	.sr_32(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[32]~q ),
	.sr_22(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[22]~q ),
	.sr_19(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[19]~q ),
	.sr_18(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[18]~q ),
	.sr_23(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[23]~q ),
	.sr_24(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[24]~q ),
	.sr_8(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[8]~q ),
	.sr_16(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[16]~q ),
	.sr_9(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[9]~q ),
	.sr_10(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[10]~q ),
	.sr_11(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[11]~q ),
	.sr_13(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[13]~q ),
	.sr_14(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[14]~q ),
	.sr_12(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[12]~q ),
	.sr_0(sr_0),
	.virtual_state_uir(\embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_uir~combout ),
	.jdo_0(jdo_0),
	.jdo_36(jdo_36),
	.jdo_37(jdo_37),
	.ir_1(ir_1),
	.ir_0(ir_0),
	.enable_action_strobe1(enable_action_strobe),
	.jdo_3(jdo_3),
	.take_action_ocimem_a1(take_action_ocimem_a),
	.jdo_35(jdo_35),
	.take_action_ocimem_b1(take_action_ocimem_b),
	.take_action_ocimem_a2(take_action_ocimem_a1),
	.jdo_34(jdo_34),
	.take_action_ocimem_a3(take_action_ocimem_a2),
	.jdo_25(jdo_25),
	.jdo_1(jdo_1),
	.jdo_4(jdo_4),
	.sr_36(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[36]~q ),
	.sr_37(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[37]~q ),
	.sr_35(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[35]~q ),
	.jdo_21(jdo_21),
	.jdo_20(jdo_20),
	.jdo_17(jdo_17),
	.sr_34(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[34]~q ),
	.jdo_2(jdo_2),
	.jdo_5(jdo_5),
	.jdo_27(jdo_27),
	.jdo_26(jdo_26),
	.jdo_28(jdo_28),
	.jdo_29(jdo_29),
	.jdo_30(jdo_30),
	.jdo_31(jdo_31),
	.jdo_32(jdo_32),
	.jdo_33(jdo_33),
	.jdo_19(jdo_19),
	.jdo_18(jdo_18),
	.jdo_6(jdo_6),
	.sr_31(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[31]~q ),
	.sr_33(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[33]~q ),
	.jdo_24(jdo_24),
	.sr_7(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[7]~q ),
	.jdo_7(jdo_7),
	.virtual_state_udr(\embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_udr~0_combout ),
	.jdo_23(jdo_23),
	.jdo_22(jdo_22),
	.jdo_16(jdo_16),
	.jdo_8(jdo_8),
	.jdo_9(jdo_9),
	.jdo_10(jdo_10),
	.jdo_15(jdo_15),
	.jdo_13(jdo_13),
	.jdo_14(jdo_14),
	.jdo_12(jdo_12),
	.jdo_11(jdo_11),
	.sr_15(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[15]~q ),
	.ir_in({irf_reg_1_1,irf_reg_0_1}),
	.clk_clk(clk_clk));

embedded_system_embedded_system_nios2_qsys_0_jtag_debug_module_tck the_embedded_system_nios2_qsys_0_jtag_debug_module_tck(
	.sr_1(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[1]~q ),
	.sr_2(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[2]~q ),
	.break_readreg_0(break_readreg_0),
	.MonDReg_0(MonDReg_0),
	.sr_3(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[3]~q ),
	.break_readreg_1(break_readreg_1),
	.sr_4(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[4]~q ),
	.break_readreg_2(break_readreg_2),
	.sr_25(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[25]~q ),
	.sr_5(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[5]~q ),
	.break_readreg_3(break_readreg_3),
	.sr_21(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[21]~q ),
	.sr_20(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[20]~q ),
	.sr_17(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[17]~q ),
	.sr_26(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[26]~q ),
	.break_readreg_24(break_readreg_24),
	.MonDReg_24(MonDReg_24),
	.sr_6(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[6]~q ),
	.break_readreg_4(break_readreg_4),
	.MonDReg_4(MonDReg_4),
	.sr_27(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[27]~q ),
	.sr_28(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[28]~q ),
	.sr_29(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[29]~q ),
	.sr_30(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[30]~q ),
	.sr_32(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[32]~q ),
	.sr_22(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[22]~q ),
	.break_readreg_20(break_readreg_20),
	.MonDReg_20(MonDReg_20),
	.break_readreg_19(break_readreg_19),
	.MonDReg_19(MonDReg_19),
	.sr_19(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[19]~q ),
	.sr_18(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[18]~q ),
	.break_readreg_16(break_readreg_16),
	.MonDReg_16(MonDReg_16),
	.break_readreg_25(break_readreg_25),
	.MonDReg_25(MonDReg_25),
	.break_readreg_5(break_readreg_5),
	.break_readreg_26(break_readreg_26),
	.MonDReg_26(MonDReg_26),
	.break_readreg_27(break_readreg_27),
	.MonDReg_27(MonDReg_27),
	.break_readreg_28(break_readreg_28),
	.MonDReg_28(MonDReg_28),
	.break_readreg_29(break_readreg_29),
	.MonDReg_30(MonDReg_30),
	.break_readreg_30(break_readreg_30),
	.break_readreg_31(break_readreg_31),
	.MonDReg_31(MonDReg_31),
	.sr_23(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[23]~q ),
	.break_readreg_21(break_readreg_21),
	.MonDReg_21(MonDReg_21),
	.break_readreg_18(break_readreg_18),
	.break_readreg_17(break_readreg_17),
	.MonDReg_17(MonDReg_17),
	.sr_24(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[24]~q ),
	.sr_8(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[8]~q ),
	.break_readreg_6(break_readreg_6),
	.MonDReg_6(MonDReg_6),
	.break_readreg_22(break_readreg_22),
	.MonDReg_22(MonDReg_22),
	.sr_16(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[16]~q ),
	.break_readreg_23(break_readreg_23),
	.MonDReg_23(MonDReg_23),
	.sr_9(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[9]~q ),
	.break_readreg_7(break_readreg_7),
	.MonDReg_7(MonDReg_7),
	.MonDReg_15(MonDReg_15),
	.break_readreg_15(break_readreg_15),
	.MonDReg_13(MonDReg_13),
	.MonDReg_14(MonDReg_14),
	.sr_10(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[10]~q ),
	.break_readreg_8(break_readreg_8),
	.sr_11(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[11]~q ),
	.break_readreg_9(break_readreg_9),
	.sr_13(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[13]~q ),
	.sr_14(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[14]~q ),
	.sr_12(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[12]~q ),
	.break_readreg_10(break_readreg_10),
	.break_readreg_14(break_readreg_14),
	.break_readreg_12(break_readreg_12),
	.break_readreg_13(break_readreg_13),
	.break_readreg_11(break_readreg_11),
	.sr_0(sr_0),
	.ir_out_0(ir_out_0),
	.ir_out_1(ir_out_1),
	.virtual_state_sdr(\embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_sdr~0_combout ),
	.virtual_state_uir(\embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_uir~combout ),
	.monitor_ready(monitor_ready),
	.MonDReg_1(MonDReg_1),
	.hbreak_enabled(hbreak_enabled),
	.MonDReg_2(MonDReg_2),
	.sr_36(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[36]~q ),
	.sr_37(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[37]~q ),
	.sr_35(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[35]~q ),
	.sr_34(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[34]~q ),
	.MonDReg_3(MonDReg_3),
	.virtual_state_cdr(\embedded_system_nios2_qsys_0_jtag_debug_module_phy|virtual_state_cdr~combout ),
	.monitor_error(monitor_error),
	.sr_31(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[31]~q ),
	.sr_33(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[33]~q ),
	.sr_7(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[7]~q ),
	.MonDReg_5(MonDReg_5),
	.MonDReg_29(MonDReg_29),
	.resetlatch(resetlatch),
	.MonDReg_18(MonDReg_18),
	.MonDReg_10(MonDReg_10),
	.MonDReg_12(MonDReg_12),
	.MonDReg_11(MonDReg_11),
	.MonDReg_9(MonDReg_9),
	.MonDReg_8(MonDReg_8),
	.sr_15(\the_embedded_system_nios2_qsys_0_jtag_debug_module_tck|sr[15]~q ),
	.altera_internal_jtag(altera_internal_jtag),
	.altera_internal_jtag1(altera_internal_jtag1),
	.state_4(state_4),
	.splitter_nodes_receive_0_3(splitter_nodes_receive_0_3),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1));

endmodule

module embedded_system_embedded_system_nios2_qsys_0_jtag_debug_module_sysclk (
	sr_1,
	sr_2,
	sr_3,
	sr_4,
	sr_25,
	sr_5,
	sr_21,
	sr_20,
	sr_17,
	sr_26,
	sr_6,
	sr_27,
	sr_28,
	sr_29,
	sr_30,
	sr_32,
	sr_22,
	sr_19,
	sr_18,
	sr_23,
	sr_24,
	sr_8,
	sr_16,
	sr_9,
	sr_10,
	sr_11,
	sr_13,
	sr_14,
	sr_12,
	sr_0,
	virtual_state_uir,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe1,
	jdo_3,
	take_action_ocimem_a1,
	jdo_35,
	take_action_ocimem_b1,
	take_action_ocimem_a2,
	jdo_34,
	take_action_ocimem_a3,
	jdo_25,
	jdo_1,
	jdo_4,
	sr_36,
	sr_37,
	sr_35,
	jdo_21,
	jdo_20,
	jdo_17,
	sr_34,
	jdo_2,
	jdo_5,
	jdo_27,
	jdo_26,
	jdo_28,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	jdo_19,
	jdo_18,
	jdo_6,
	sr_31,
	sr_33,
	jdo_24,
	sr_7,
	jdo_7,
	virtual_state_udr,
	jdo_23,
	jdo_22,
	jdo_16,
	jdo_8,
	jdo_9,
	jdo_10,
	jdo_15,
	jdo_13,
	jdo_14,
	jdo_12,
	jdo_11,
	sr_15,
	ir_in,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	sr_1;
input 	sr_2;
input 	sr_3;
input 	sr_4;
input 	sr_25;
input 	sr_5;
input 	sr_21;
input 	sr_20;
input 	sr_17;
input 	sr_26;
input 	sr_6;
input 	sr_27;
input 	sr_28;
input 	sr_29;
input 	sr_30;
input 	sr_32;
input 	sr_22;
input 	sr_19;
input 	sr_18;
input 	sr_23;
input 	sr_24;
input 	sr_8;
input 	sr_16;
input 	sr_9;
input 	sr_10;
input 	sr_11;
input 	sr_13;
input 	sr_14;
input 	sr_12;
input 	sr_0;
input 	virtual_state_uir;
output 	jdo_0;
output 	jdo_36;
output 	jdo_37;
output 	ir_1;
output 	ir_0;
output 	enable_action_strobe1;
output 	jdo_3;
output 	take_action_ocimem_a1;
output 	jdo_35;
output 	take_action_ocimem_b1;
output 	take_action_ocimem_a2;
output 	jdo_34;
output 	take_action_ocimem_a3;
output 	jdo_25;
output 	jdo_1;
output 	jdo_4;
input 	sr_36;
input 	sr_37;
input 	sr_35;
output 	jdo_21;
output 	jdo_20;
output 	jdo_17;
input 	sr_34;
output 	jdo_2;
output 	jdo_5;
output 	jdo_27;
output 	jdo_26;
output 	jdo_28;
output 	jdo_29;
output 	jdo_30;
output 	jdo_31;
output 	jdo_32;
output 	jdo_33;
output 	jdo_19;
output 	jdo_18;
output 	jdo_6;
input 	sr_31;
input 	sr_33;
output 	jdo_24;
input 	sr_7;
output 	jdo_7;
input 	virtual_state_udr;
output 	jdo_23;
output 	jdo_22;
output 	jdo_16;
output 	jdo_8;
output 	jdo_9;
output 	jdo_10;
output 	jdo_15;
output 	jdo_13;
output 	jdo_14;
output 	jdo_12;
output 	jdo_11;
input 	sr_15;
input 	[1:0] ir_in;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer3|dreg[0]~q ;
wire \the_altera_std_synchronizer4|dreg[0]~q ;
wire \sync2_udr~q ;
wire \update_jdo_strobe~0_combout ;
wire \update_jdo_strobe~q ;
wire \sync2_uir~q ;
wire \jxuir~0_combout ;
wire \jxuir~q ;


embedded_system_altera_std_synchronizer_1 the_altera_std_synchronizer4(
	.din(virtual_state_uir),
	.dreg_0(\the_altera_std_synchronizer4|dreg[0]~q ),
	.clk(clk_clk));

embedded_system_altera_std_synchronizer the_altera_std_synchronizer3(
	.dreg_0(\the_altera_std_synchronizer3|dreg[0]~q ),
	.din(virtual_state_udr),
	.clk(clk_clk));

dffeas \jdo[0] (
	.clk(clk_clk),
	.d(sr_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_0),
	.prn(vcc));
defparam \jdo[0] .is_wysiwyg = "true";
defparam \jdo[0] .power_up = "low";

dffeas \jdo[36] (
	.clk(clk_clk),
	.d(sr_36),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_36),
	.prn(vcc));
defparam \jdo[36] .is_wysiwyg = "true";
defparam \jdo[36] .power_up = "low";

dffeas \jdo[37] (
	.clk(clk_clk),
	.d(sr_37),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_37),
	.prn(vcc));
defparam \jdo[37] .is_wysiwyg = "true";
defparam \jdo[37] .power_up = "low";

dffeas \ir[1] (
	.clk(clk_clk),
	.d(ir_in[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_1),
	.prn(vcc));
defparam \ir[1] .is_wysiwyg = "true";
defparam \ir[1] .power_up = "low";

dffeas \ir[0] (
	.clk(clk_clk),
	.d(ir_in[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\jxuir~q ),
	.q(ir_0),
	.prn(vcc));
defparam \ir[0] .is_wysiwyg = "true";
defparam \ir[0] .power_up = "low";

dffeas enable_action_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(enable_action_strobe1),
	.prn(vcc));
defparam enable_action_strobe.is_wysiwyg = "true";
defparam enable_action_strobe.power_up = "low";

dffeas \jdo[3] (
	.clk(clk_clk),
	.d(sr_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_3),
	.prn(vcc));
defparam \jdo[3] .is_wysiwyg = "true";
defparam \jdo[3] .power_up = "low";

cyclonev_lcell_comb \take_action_ocimem_a~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a1),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~0 .extended_lut = "off";
defparam \take_action_ocimem_a~0 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \take_action_ocimem_a~0 .shared_arith = "off";

dffeas \jdo[35] (
	.clk(clk_clk),
	.d(sr_35),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_35),
	.prn(vcc));
defparam \jdo[35] .is_wysiwyg = "true";
defparam \jdo[35] .power_up = "low";

cyclonev_lcell_comb take_action_ocimem_b(
	.dataa(!take_action_ocimem_a1),
	.datab(!jdo_35),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_b1),
	.sumout(),
	.cout(),
	.shareout());
defparam take_action_ocimem_b.extended_lut = "off";
defparam take_action_ocimem_b.lut_mask = 64'h7777777777777777;
defparam take_action_ocimem_b.shared_arith = "off";

cyclonev_lcell_comb \take_action_ocimem_a~1 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe1),
	.datad(!jdo_35),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a2),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocimem_a~1 .extended_lut = "off";
defparam \take_action_ocimem_a~1 .lut_mask = 64'hFFEFFFEFFFEFFFEF;
defparam \take_action_ocimem_a~1 .shared_arith = "off";

dffeas \jdo[34] (
	.clk(clk_clk),
	.d(sr_34),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_34),
	.prn(vcc));
defparam \jdo[34] .is_wysiwyg = "true";
defparam \jdo[34] .power_up = "low";

cyclonev_lcell_comb take_action_ocimem_a(
	.dataa(!take_action_ocimem_a2),
	.datab(!jdo_34),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocimem_a3),
	.sumout(),
	.cout(),
	.shareout());
defparam take_action_ocimem_a.extended_lut = "off";
defparam take_action_ocimem_a.lut_mask = 64'h7777777777777777;
defparam take_action_ocimem_a.shared_arith = "off";

dffeas \jdo[25] (
	.clk(clk_clk),
	.d(sr_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_25),
	.prn(vcc));
defparam \jdo[25] .is_wysiwyg = "true";
defparam \jdo[25] .power_up = "low";

dffeas \jdo[1] (
	.clk(clk_clk),
	.d(sr_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_1),
	.prn(vcc));
defparam \jdo[1] .is_wysiwyg = "true";
defparam \jdo[1] .power_up = "low";

dffeas \jdo[4] (
	.clk(clk_clk),
	.d(sr_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_4),
	.prn(vcc));
defparam \jdo[4] .is_wysiwyg = "true";
defparam \jdo[4] .power_up = "low";

dffeas \jdo[21] (
	.clk(clk_clk),
	.d(sr_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_21),
	.prn(vcc));
defparam \jdo[21] .is_wysiwyg = "true";
defparam \jdo[21] .power_up = "low";

dffeas \jdo[20] (
	.clk(clk_clk),
	.d(sr_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_20),
	.prn(vcc));
defparam \jdo[20] .is_wysiwyg = "true";
defparam \jdo[20] .power_up = "low";

dffeas \jdo[17] (
	.clk(clk_clk),
	.d(sr_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_17),
	.prn(vcc));
defparam \jdo[17] .is_wysiwyg = "true";
defparam \jdo[17] .power_up = "low";

dffeas \jdo[2] (
	.clk(clk_clk),
	.d(sr_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_2),
	.prn(vcc));
defparam \jdo[2] .is_wysiwyg = "true";
defparam \jdo[2] .power_up = "low";

dffeas \jdo[5] (
	.clk(clk_clk),
	.d(sr_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_5),
	.prn(vcc));
defparam \jdo[5] .is_wysiwyg = "true";
defparam \jdo[5] .power_up = "low";

dffeas \jdo[27] (
	.clk(clk_clk),
	.d(sr_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_27),
	.prn(vcc));
defparam \jdo[27] .is_wysiwyg = "true";
defparam \jdo[27] .power_up = "low";

dffeas \jdo[26] (
	.clk(clk_clk),
	.d(sr_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_26),
	.prn(vcc));
defparam \jdo[26] .is_wysiwyg = "true";
defparam \jdo[26] .power_up = "low";

dffeas \jdo[28] (
	.clk(clk_clk),
	.d(sr_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_28),
	.prn(vcc));
defparam \jdo[28] .is_wysiwyg = "true";
defparam \jdo[28] .power_up = "low";

dffeas \jdo[29] (
	.clk(clk_clk),
	.d(sr_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_29),
	.prn(vcc));
defparam \jdo[29] .is_wysiwyg = "true";
defparam \jdo[29] .power_up = "low";

dffeas \jdo[30] (
	.clk(clk_clk),
	.d(sr_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_30),
	.prn(vcc));
defparam \jdo[30] .is_wysiwyg = "true";
defparam \jdo[30] .power_up = "low";

dffeas \jdo[31] (
	.clk(clk_clk),
	.d(sr_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_31),
	.prn(vcc));
defparam \jdo[31] .is_wysiwyg = "true";
defparam \jdo[31] .power_up = "low";

dffeas \jdo[32] (
	.clk(clk_clk),
	.d(sr_32),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_32),
	.prn(vcc));
defparam \jdo[32] .is_wysiwyg = "true";
defparam \jdo[32] .power_up = "low";

dffeas \jdo[33] (
	.clk(clk_clk),
	.d(sr_33),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_33),
	.prn(vcc));
defparam \jdo[33] .is_wysiwyg = "true";
defparam \jdo[33] .power_up = "low";

dffeas \jdo[19] (
	.clk(clk_clk),
	.d(sr_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_19),
	.prn(vcc));
defparam \jdo[19] .is_wysiwyg = "true";
defparam \jdo[19] .power_up = "low";

dffeas \jdo[18] (
	.clk(clk_clk),
	.d(sr_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_18),
	.prn(vcc));
defparam \jdo[18] .is_wysiwyg = "true";
defparam \jdo[18] .power_up = "low";

dffeas \jdo[6] (
	.clk(clk_clk),
	.d(sr_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_6),
	.prn(vcc));
defparam \jdo[6] .is_wysiwyg = "true";
defparam \jdo[6] .power_up = "low";

dffeas \jdo[24] (
	.clk(clk_clk),
	.d(sr_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_24),
	.prn(vcc));
defparam \jdo[24] .is_wysiwyg = "true";
defparam \jdo[24] .power_up = "low";

dffeas \jdo[7] (
	.clk(clk_clk),
	.d(sr_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_7),
	.prn(vcc));
defparam \jdo[7] .is_wysiwyg = "true";
defparam \jdo[7] .power_up = "low";

dffeas \jdo[23] (
	.clk(clk_clk),
	.d(sr_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_23),
	.prn(vcc));
defparam \jdo[23] .is_wysiwyg = "true";
defparam \jdo[23] .power_up = "low";

dffeas \jdo[22] (
	.clk(clk_clk),
	.d(sr_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_22),
	.prn(vcc));
defparam \jdo[22] .is_wysiwyg = "true";
defparam \jdo[22] .power_up = "low";

dffeas \jdo[16] (
	.clk(clk_clk),
	.d(sr_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_16),
	.prn(vcc));
defparam \jdo[16] .is_wysiwyg = "true";
defparam \jdo[16] .power_up = "low";

dffeas \jdo[8] (
	.clk(clk_clk),
	.d(sr_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_8),
	.prn(vcc));
defparam \jdo[8] .is_wysiwyg = "true";
defparam \jdo[8] .power_up = "low";

dffeas \jdo[9] (
	.clk(clk_clk),
	.d(sr_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_9),
	.prn(vcc));
defparam \jdo[9] .is_wysiwyg = "true";
defparam \jdo[9] .power_up = "low";

dffeas \jdo[10] (
	.clk(clk_clk),
	.d(sr_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_10),
	.prn(vcc));
defparam \jdo[10] .is_wysiwyg = "true";
defparam \jdo[10] .power_up = "low";

dffeas \jdo[15] (
	.clk(clk_clk),
	.d(sr_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_15),
	.prn(vcc));
defparam \jdo[15] .is_wysiwyg = "true";
defparam \jdo[15] .power_up = "low";

dffeas \jdo[13] (
	.clk(clk_clk),
	.d(sr_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_13),
	.prn(vcc));
defparam \jdo[13] .is_wysiwyg = "true";
defparam \jdo[13] .power_up = "low";

dffeas \jdo[14] (
	.clk(clk_clk),
	.d(sr_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_14),
	.prn(vcc));
defparam \jdo[14] .is_wysiwyg = "true";
defparam \jdo[14] .power_up = "low";

dffeas \jdo[12] (
	.clk(clk_clk),
	.d(sr_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_12),
	.prn(vcc));
defparam \jdo[12] .is_wysiwyg = "true";
defparam \jdo[12] .power_up = "low";

dffeas \jdo[11] (
	.clk(clk_clk),
	.d(sr_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\update_jdo_strobe~q ),
	.q(jdo_11),
	.prn(vcc));
defparam \jdo[11] .is_wysiwyg = "true";
defparam \jdo[11] .power_up = "low";

dffeas sync2_udr(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer3|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_udr~q ),
	.prn(vcc));
defparam sync2_udr.is_wysiwyg = "true";
defparam sync2_udr.power_up = "low";

cyclonev_lcell_comb \update_jdo_strobe~0 (
	.dataa(!\sync2_udr~q ),
	.datab(!\the_altera_std_synchronizer3|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\update_jdo_strobe~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \update_jdo_strobe~0 .extended_lut = "off";
defparam \update_jdo_strobe~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \update_jdo_strobe~0 .shared_arith = "off";

dffeas update_jdo_strobe(
	.clk(clk_clk),
	.d(\update_jdo_strobe~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\update_jdo_strobe~q ),
	.prn(vcc));
defparam update_jdo_strobe.is_wysiwyg = "true";
defparam update_jdo_strobe.power_up = "low";

dffeas sync2_uir(
	.clk(clk_clk),
	.d(\the_altera_std_synchronizer4|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sync2_uir~q ),
	.prn(vcc));
defparam sync2_uir.is_wysiwyg = "true";
defparam sync2_uir.power_up = "low";

cyclonev_lcell_comb \jxuir~0 (
	.dataa(!\sync2_uir~q ),
	.datab(!\the_altera_std_synchronizer4|dreg[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jxuir~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jxuir~0 .extended_lut = "off";
defparam \jxuir~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \jxuir~0 .shared_arith = "off";

dffeas jxuir(
	.clk(clk_clk),
	.d(\jxuir~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jxuir~q ),
	.prn(vcc));
defparam jxuir.is_wysiwyg = "true";
defparam jxuir.power_up = "low";

endmodule

module embedded_system_altera_std_synchronizer (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module embedded_system_altera_std_synchronizer_1 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_jtag_debug_module_tck (
	sr_1,
	sr_2,
	break_readreg_0,
	MonDReg_0,
	sr_3,
	break_readreg_1,
	sr_4,
	break_readreg_2,
	sr_25,
	sr_5,
	break_readreg_3,
	sr_21,
	sr_20,
	sr_17,
	sr_26,
	break_readreg_24,
	MonDReg_24,
	sr_6,
	break_readreg_4,
	MonDReg_4,
	sr_27,
	sr_28,
	sr_29,
	sr_30,
	sr_32,
	sr_22,
	break_readreg_20,
	MonDReg_20,
	break_readreg_19,
	MonDReg_19,
	sr_19,
	sr_18,
	break_readreg_16,
	MonDReg_16,
	break_readreg_25,
	MonDReg_25,
	break_readreg_5,
	break_readreg_26,
	MonDReg_26,
	break_readreg_27,
	MonDReg_27,
	break_readreg_28,
	MonDReg_28,
	break_readreg_29,
	MonDReg_30,
	break_readreg_30,
	break_readreg_31,
	MonDReg_31,
	sr_23,
	break_readreg_21,
	MonDReg_21,
	break_readreg_18,
	break_readreg_17,
	MonDReg_17,
	sr_24,
	sr_8,
	break_readreg_6,
	MonDReg_6,
	break_readreg_22,
	MonDReg_22,
	sr_16,
	break_readreg_23,
	MonDReg_23,
	sr_9,
	break_readreg_7,
	MonDReg_7,
	MonDReg_15,
	break_readreg_15,
	MonDReg_13,
	MonDReg_14,
	sr_10,
	break_readreg_8,
	sr_11,
	break_readreg_9,
	sr_13,
	sr_14,
	sr_12,
	break_readreg_10,
	break_readreg_14,
	break_readreg_12,
	break_readreg_13,
	break_readreg_11,
	sr_0,
	ir_out_0,
	ir_out_1,
	virtual_state_sdr,
	virtual_state_uir,
	monitor_ready,
	MonDReg_1,
	hbreak_enabled,
	MonDReg_2,
	sr_36,
	sr_37,
	sr_35,
	sr_34,
	MonDReg_3,
	virtual_state_cdr,
	monitor_error,
	sr_31,
	sr_33,
	sr_7,
	MonDReg_5,
	MonDReg_29,
	resetlatch,
	MonDReg_18,
	MonDReg_10,
	MonDReg_12,
	MonDReg_11,
	MonDReg_9,
	MonDReg_8,
	sr_15,
	altera_internal_jtag,
	altera_internal_jtag1,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	irf_reg_0_1,
	irf_reg_1_1)/* synthesis synthesis_greybox=1 */;
output 	sr_1;
output 	sr_2;
input 	break_readreg_0;
input 	MonDReg_0;
output 	sr_3;
input 	break_readreg_1;
output 	sr_4;
input 	break_readreg_2;
output 	sr_25;
output 	sr_5;
input 	break_readreg_3;
output 	sr_21;
output 	sr_20;
output 	sr_17;
output 	sr_26;
input 	break_readreg_24;
input 	MonDReg_24;
output 	sr_6;
input 	break_readreg_4;
input 	MonDReg_4;
output 	sr_27;
output 	sr_28;
output 	sr_29;
output 	sr_30;
output 	sr_32;
output 	sr_22;
input 	break_readreg_20;
input 	MonDReg_20;
input 	break_readreg_19;
input 	MonDReg_19;
output 	sr_19;
output 	sr_18;
input 	break_readreg_16;
input 	MonDReg_16;
input 	break_readreg_25;
input 	MonDReg_25;
input 	break_readreg_5;
input 	break_readreg_26;
input 	MonDReg_26;
input 	break_readreg_27;
input 	MonDReg_27;
input 	break_readreg_28;
input 	MonDReg_28;
input 	break_readreg_29;
input 	MonDReg_30;
input 	break_readreg_30;
input 	break_readreg_31;
input 	MonDReg_31;
output 	sr_23;
input 	break_readreg_21;
input 	MonDReg_21;
input 	break_readreg_18;
input 	break_readreg_17;
input 	MonDReg_17;
output 	sr_24;
output 	sr_8;
input 	break_readreg_6;
input 	MonDReg_6;
input 	break_readreg_22;
input 	MonDReg_22;
output 	sr_16;
input 	break_readreg_23;
input 	MonDReg_23;
output 	sr_9;
input 	break_readreg_7;
input 	MonDReg_7;
input 	MonDReg_15;
input 	break_readreg_15;
input 	MonDReg_13;
input 	MonDReg_14;
output 	sr_10;
input 	break_readreg_8;
output 	sr_11;
input 	break_readreg_9;
output 	sr_13;
output 	sr_14;
output 	sr_12;
input 	break_readreg_10;
input 	break_readreg_14;
input 	break_readreg_12;
input 	break_readreg_13;
input 	break_readreg_11;
output 	sr_0;
output 	ir_out_0;
output 	ir_out_1;
input 	virtual_state_sdr;
input 	virtual_state_uir;
input 	monitor_ready;
input 	MonDReg_1;
input 	hbreak_enabled;
input 	MonDReg_2;
output 	sr_36;
output 	sr_37;
output 	sr_35;
output 	sr_34;
input 	MonDReg_3;
input 	virtual_state_cdr;
input 	monitor_error;
output 	sr_31;
output 	sr_33;
output 	sr_7;
input 	MonDReg_5;
input 	MonDReg_29;
input 	resetlatch;
input 	MonDReg_18;
input 	MonDReg_10;
input 	MonDReg_12;
input 	MonDReg_11;
input 	MonDReg_9;
input 	MonDReg_8;
output 	sr_15;
input 	altera_internal_jtag;
input 	altera_internal_jtag1;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	irf_reg_0_1;
input 	irf_reg_1_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer2|dreg[0]~q ;
wire \the_altera_std_synchronizer1|dreg[0]~q ;
wire \sr~8_combout ;
wire \sr[2]~9_combout ;
wire \sr[2]~10_combout ;
wire \sr~11_combout ;
wire \sr~12_combout ;
wire \sr~13_combout ;
wire \sr~20_combout ;
wire \sr[23]~21_combout ;
wire \sr[23]~19_combout ;
wire \sr~22_combout ;
wire \sr~23_combout ;
wire \sr~24_combout ;
wire \sr~25_combout ;
wire \sr~26_combout ;
wire \sr~27_combout ;
wire \sr~28_combout ;
wire \sr~29_combout ;
wire \sr~30_combout ;
wire \sr~31_combout ;
wire \sr~36_combout ;
wire \sr~38_combout ;
wire \sr~39_combout ;
wire \sr~40_combout ;
wire \sr~43_combout ;
wire \sr~44_combout ;
wire \sr~45_combout ;
wire \sr~46_combout ;
wire \sr~47_combout ;
wire \sr~48_combout ;
wire \sr~49_combout ;
wire \sr~52_combout ;
wire \sr~53_combout ;
wire \sr~54_combout ;
wire \sr~5_combout ;
wire \sr~6_combout ;
wire \DRsize.000~q ;
wire \sr~7_combout ;
wire \sr~14_combout ;
wire \sr[36]~15_combout ;
wire \sr~16_combout ;
wire \Mux37~0_combout ;
wire \DRsize.100~q ;
wire \sr~56_combout ;
wire \sr~17_combout ;
wire \sr~18_combout ;
wire \sr[23]~32_combout ;
wire \sr~33_combout ;
wire \sr~34_combout ;
wire \sr~35_combout ;
wire \sr~37_combout ;
wire \sr~41_combout ;
wire \sr~42_combout ;
wire \sr[23]~55_combout ;
wire \DRsize.010~q ;
wire \sr~50_combout ;
wire \sr~51_combout ;


embedded_system_altera_std_synchronizer_3 the_altera_std_synchronizer2(
	.dreg_0(\the_altera_std_synchronizer2|dreg[0]~q ),
	.din(monitor_ready),
	.clk(altera_internal_jtag));

embedded_system_altera_std_synchronizer_2 the_altera_std_synchronizer1(
	.dreg_0(\the_altera_std_synchronizer1|dreg[0]~q ),
	.din(hbreak_enabled),
	.clk(altera_internal_jtag));

dffeas \sr[1] (
	.clk(altera_internal_jtag),
	.d(\sr~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_1),
	.prn(vcc));
defparam \sr[1] .is_wysiwyg = "true";
defparam \sr[1] .power_up = "low";

dffeas \sr[2] (
	.clk(altera_internal_jtag),
	.d(\sr~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_2),
	.prn(vcc));
defparam \sr[2] .is_wysiwyg = "true";
defparam \sr[2] .power_up = "low";

dffeas \sr[3] (
	.clk(altera_internal_jtag),
	.d(\sr~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_3),
	.prn(vcc));
defparam \sr[3] .is_wysiwyg = "true";
defparam \sr[3] .power_up = "low";

dffeas \sr[4] (
	.clk(altera_internal_jtag),
	.d(\sr~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_4),
	.prn(vcc));
defparam \sr[4] .is_wysiwyg = "true";
defparam \sr[4] .power_up = "low";

dffeas \sr[25] (
	.clk(altera_internal_jtag),
	.d(\sr~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_25),
	.prn(vcc));
defparam \sr[25] .is_wysiwyg = "true";
defparam \sr[25] .power_up = "low";

dffeas \sr[5] (
	.clk(altera_internal_jtag),
	.d(\sr~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_5),
	.prn(vcc));
defparam \sr[5] .is_wysiwyg = "true";
defparam \sr[5] .power_up = "low";

dffeas \sr[21] (
	.clk(altera_internal_jtag),
	.d(\sr~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_21),
	.prn(vcc));
defparam \sr[21] .is_wysiwyg = "true";
defparam \sr[21] .power_up = "low";

dffeas \sr[20] (
	.clk(altera_internal_jtag),
	.d(\sr~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_20),
	.prn(vcc));
defparam \sr[20] .is_wysiwyg = "true";
defparam \sr[20] .power_up = "low";

dffeas \sr[17] (
	.clk(altera_internal_jtag),
	.d(\sr~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_17),
	.prn(vcc));
defparam \sr[17] .is_wysiwyg = "true";
defparam \sr[17] .power_up = "low";

dffeas \sr[26] (
	.clk(altera_internal_jtag),
	.d(\sr~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_26),
	.prn(vcc));
defparam \sr[26] .is_wysiwyg = "true";
defparam \sr[26] .power_up = "low";

dffeas \sr[6] (
	.clk(altera_internal_jtag),
	.d(\sr~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_6),
	.prn(vcc));
defparam \sr[6] .is_wysiwyg = "true";
defparam \sr[6] .power_up = "low";

dffeas \sr[27] (
	.clk(altera_internal_jtag),
	.d(\sr~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_27),
	.prn(vcc));
defparam \sr[27] .is_wysiwyg = "true";
defparam \sr[27] .power_up = "low";

dffeas \sr[28] (
	.clk(altera_internal_jtag),
	.d(\sr~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_28),
	.prn(vcc));
defparam \sr[28] .is_wysiwyg = "true";
defparam \sr[28] .power_up = "low";

dffeas \sr[29] (
	.clk(altera_internal_jtag),
	.d(\sr~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_29),
	.prn(vcc));
defparam \sr[29] .is_wysiwyg = "true";
defparam \sr[29] .power_up = "low";

dffeas \sr[30] (
	.clk(altera_internal_jtag),
	.d(\sr~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_30),
	.prn(vcc));
defparam \sr[30] .is_wysiwyg = "true";
defparam \sr[30] .power_up = "low";

dffeas \sr[32] (
	.clk(altera_internal_jtag),
	.d(\sr~36_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_32),
	.prn(vcc));
defparam \sr[32] .is_wysiwyg = "true";
defparam \sr[32] .power_up = "low";

dffeas \sr[22] (
	.clk(altera_internal_jtag),
	.d(\sr~38_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_22),
	.prn(vcc));
defparam \sr[22] .is_wysiwyg = "true";
defparam \sr[22] .power_up = "low";

dffeas \sr[19] (
	.clk(altera_internal_jtag),
	.d(\sr~39_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_19),
	.prn(vcc));
defparam \sr[19] .is_wysiwyg = "true";
defparam \sr[19] .power_up = "low";

dffeas \sr[18] (
	.clk(altera_internal_jtag),
	.d(\sr~40_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_18),
	.prn(vcc));
defparam \sr[18] .is_wysiwyg = "true";
defparam \sr[18] .power_up = "low";

dffeas \sr[23] (
	.clk(altera_internal_jtag),
	.d(\sr~43_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_23),
	.prn(vcc));
defparam \sr[23] .is_wysiwyg = "true";
defparam \sr[23] .power_up = "low";

dffeas \sr[24] (
	.clk(altera_internal_jtag),
	.d(\sr~44_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_24),
	.prn(vcc));
defparam \sr[24] .is_wysiwyg = "true";
defparam \sr[24] .power_up = "low";

dffeas \sr[8] (
	.clk(altera_internal_jtag),
	.d(\sr~45_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_8),
	.prn(vcc));
defparam \sr[8] .is_wysiwyg = "true";
defparam \sr[8] .power_up = "low";

dffeas \sr[16] (
	.clk(altera_internal_jtag),
	.d(\sr~46_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[23]~21_combout ),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_16),
	.prn(vcc));
defparam \sr[16] .is_wysiwyg = "true";
defparam \sr[16] .power_up = "low";

dffeas \sr[9] (
	.clk(altera_internal_jtag),
	.d(\sr~47_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_9),
	.prn(vcc));
defparam \sr[9] .is_wysiwyg = "true";
defparam \sr[9] .power_up = "low";

dffeas \sr[10] (
	.clk(altera_internal_jtag),
	.d(\sr~48_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_10),
	.prn(vcc));
defparam \sr[10] .is_wysiwyg = "true";
defparam \sr[10] .power_up = "low";

dffeas \sr[11] (
	.clk(altera_internal_jtag),
	.d(\sr~49_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_11),
	.prn(vcc));
defparam \sr[11] .is_wysiwyg = "true";
defparam \sr[11] .power_up = "low";

dffeas \sr[13] (
	.clk(altera_internal_jtag),
	.d(\sr~52_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_13),
	.prn(vcc));
defparam \sr[13] .is_wysiwyg = "true";
defparam \sr[13] .power_up = "low";

dffeas \sr[14] (
	.clk(altera_internal_jtag),
	.d(\sr~53_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_14),
	.prn(vcc));
defparam \sr[14] .is_wysiwyg = "true";
defparam \sr[14] .power_up = "low";

dffeas \sr[12] (
	.clk(altera_internal_jtag),
	.d(\sr~54_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\sr[2]~9_combout ),
	.sload(gnd),
	.ena(\sr[2]~10_combout ),
	.q(sr_12),
	.prn(vcc));
defparam \sr[12] .is_wysiwyg = "true";
defparam \sr[12] .power_up = "low";

dffeas \sr[0] (
	.clk(altera_internal_jtag),
	.d(\sr~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_0),
	.prn(vcc));
defparam \sr[0] .is_wysiwyg = "true";
defparam \sr[0] .power_up = "low";

dffeas \ir_out[0] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer2|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_0),
	.prn(vcc));
defparam \ir_out[0] .is_wysiwyg = "true";
defparam \ir_out[0] .power_up = "low";

dffeas \ir_out[1] (
	.clk(altera_internal_jtag),
	.d(\the_altera_std_synchronizer1|dreg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(ir_out_1),
	.prn(vcc));
defparam \ir_out[1] .is_wysiwyg = "true";
defparam \ir_out[1] .power_up = "low";

dffeas \sr[36] (
	.clk(altera_internal_jtag),
	.d(\sr~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[36]~15_combout ),
	.q(sr_36),
	.prn(vcc));
defparam \sr[36] .is_wysiwyg = "true";
defparam \sr[36] .power_up = "low";

dffeas \sr[37] (
	.clk(altera_internal_jtag),
	.d(\sr~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[36]~15_combout ),
	.q(sr_37),
	.prn(vcc));
defparam \sr[37] .is_wysiwyg = "true";
defparam \sr[37] .power_up = "low";

dffeas \sr[35] (
	.clk(altera_internal_jtag),
	.d(\sr~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_35),
	.prn(vcc));
defparam \sr[35] .is_wysiwyg = "true";
defparam \sr[35] .power_up = "low";

dffeas \sr[34] (
	.clk(altera_internal_jtag),
	.d(\sr~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_34),
	.prn(vcc));
defparam \sr[34] .is_wysiwyg = "true";
defparam \sr[34] .power_up = "low";

dffeas \sr[31] (
	.clk(altera_internal_jtag),
	.d(\sr~35_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_31),
	.prn(vcc));
defparam \sr[31] .is_wysiwyg = "true";
defparam \sr[31] .power_up = "low";

dffeas \sr[33] (
	.clk(altera_internal_jtag),
	.d(\sr~37_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\sr[23]~19_combout ),
	.q(sr_33),
	.prn(vcc));
defparam \sr[33] .is_wysiwyg = "true";
defparam \sr[33] .power_up = "low";

dffeas \sr[7] (
	.clk(altera_internal_jtag),
	.d(\sr~42_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_7),
	.prn(vcc));
defparam \sr[7] .is_wysiwyg = "true";
defparam \sr[7] .power_up = "low";

dffeas \sr[15] (
	.clk(altera_internal_jtag),
	.d(\sr~51_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(sr_15),
	.prn(vcc));
defparam \sr[15] .is_wysiwyg = "true";
defparam \sr[15] .power_up = "low";

cyclonev_lcell_comb \sr~8 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_2),
	.datad(!break_readreg_0),
	.datae(!MonDReg_0),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~8 .extended_lut = "off";
defparam \sr~8 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~8 .shared_arith = "off";

cyclonev_lcell_comb \sr[2]~9 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!irf_reg_0_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[2]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[2]~9 .extended_lut = "off";
defparam \sr[2]~9 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \sr[2]~9 .shared_arith = "off";

cyclonev_lcell_comb \sr[2]~10 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[2]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[2]~10 .extended_lut = "off";
defparam \sr[2]~10 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr[2]~10 .shared_arith = "off";

cyclonev_lcell_comb \sr~11 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_3),
	.datad(!break_readreg_1),
	.datae(!MonDReg_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~11 .extended_lut = "off";
defparam \sr~11 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~11 .shared_arith = "off";

cyclonev_lcell_comb \sr~12 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_4),
	.datad(!break_readreg_2),
	.datae(!MonDReg_2),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~12 .extended_lut = "off";
defparam \sr~12 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~12 .shared_arith = "off";

cyclonev_lcell_comb \sr~13 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_5),
	.datad(!break_readreg_3),
	.datae(!MonDReg_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~13 .extended_lut = "off";
defparam \sr~13 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~13 .shared_arith = "off";

cyclonev_lcell_comb \sr~20 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_26),
	.datad(!break_readreg_24),
	.datae(!MonDReg_24),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~20 .extended_lut = "off";
defparam \sr~20 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~20 .shared_arith = "off";

cyclonev_lcell_comb \sr[23]~21 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!irf_reg_0_1),
	.datae(!irf_reg_1_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[23]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[23]~21 .extended_lut = "off";
defparam \sr[23]~21 .lut_mask = 64'hFFFFFBFFFFFFFBFF;
defparam \sr[23]~21 .shared_arith = "off";

cyclonev_lcell_comb \sr[23]~19 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!state_3),
	.datae(!irf_reg_0_1),
	.dataf(!irf_reg_1_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[23]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[23]~19 .extended_lut = "off";
defparam \sr[23]~19 .lut_mask = 64'hFFFFFFFFFFFFDFFF;
defparam \sr[23]~19 .shared_arith = "off";

cyclonev_lcell_comb \sr~22 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_6),
	.datad(!break_readreg_4),
	.datae(!MonDReg_4),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~22 .extended_lut = "off";
defparam \sr~22 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~22 .shared_arith = "off";

cyclonev_lcell_comb \sr~23 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_22),
	.datad(!break_readreg_20),
	.datae(!MonDReg_20),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~23 .extended_lut = "off";
defparam \sr~23 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~23 .shared_arith = "off";

cyclonev_lcell_comb \sr~24 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_21),
	.datad(!break_readreg_19),
	.datae(!MonDReg_19),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~24 .extended_lut = "off";
defparam \sr~24 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~24 .shared_arith = "off";

cyclonev_lcell_comb \sr~25 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_18),
	.datad(!break_readreg_16),
	.datae(!MonDReg_16),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~25 .extended_lut = "off";
defparam \sr~25 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~25 .shared_arith = "off";

cyclonev_lcell_comb \sr~26 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_27),
	.datad(!break_readreg_25),
	.datae(!MonDReg_25),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~26 .extended_lut = "off";
defparam \sr~26 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~26 .shared_arith = "off";

cyclonev_lcell_comb \sr~27 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_7),
	.datad(!break_readreg_5),
	.datae(!MonDReg_5),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~27 .extended_lut = "off";
defparam \sr~27 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~27 .shared_arith = "off";

cyclonev_lcell_comb \sr~28 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_28),
	.datad(!break_readreg_26),
	.datae(!MonDReg_26),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~28 .extended_lut = "off";
defparam \sr~28 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~28 .shared_arith = "off";

cyclonev_lcell_comb \sr~29 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_29),
	.datad(!break_readreg_27),
	.datae(!MonDReg_27),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~29 .extended_lut = "off";
defparam \sr~29 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~29 .shared_arith = "off";

cyclonev_lcell_comb \sr~30 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_30),
	.datad(!break_readreg_28),
	.datae(!MonDReg_28),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~30 .extended_lut = "off";
defparam \sr~30 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~30 .shared_arith = "off";

cyclonev_lcell_comb \sr~31 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_31),
	.datad(!break_readreg_29),
	.datae(!MonDReg_29),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~31 .extended_lut = "off";
defparam \sr~31 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~31 .shared_arith = "off";

cyclonev_lcell_comb \sr~36 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_33),
	.datad(!break_readreg_31),
	.datae(!MonDReg_31),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~36_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~36 .extended_lut = "off";
defparam \sr~36 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~36 .shared_arith = "off";

cyclonev_lcell_comb \sr~38 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_23),
	.datad(!break_readreg_21),
	.datae(!MonDReg_21),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~38_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~38 .extended_lut = "off";
defparam \sr~38 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~38 .shared_arith = "off";

cyclonev_lcell_comb \sr~39 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_20),
	.datad(!break_readreg_18),
	.datae(!MonDReg_18),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~39_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~39 .extended_lut = "off";
defparam \sr~39 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~39 .shared_arith = "off";

cyclonev_lcell_comb \sr~40 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_19),
	.datad(!break_readreg_17),
	.datae(!MonDReg_17),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~40_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~40 .extended_lut = "off";
defparam \sr~40 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~40 .shared_arith = "off";

cyclonev_lcell_comb \sr~43 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_24),
	.datad(!break_readreg_22),
	.datae(!MonDReg_22),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~43_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~43 .extended_lut = "off";
defparam \sr~43 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~43 .shared_arith = "off";

cyclonev_lcell_comb \sr~44 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_25),
	.datad(!break_readreg_23),
	.datae(!MonDReg_23),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~44_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~44 .extended_lut = "off";
defparam \sr~44 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~44 .shared_arith = "off";

cyclonev_lcell_comb \sr~45 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_9),
	.datad(!break_readreg_7),
	.datae(!MonDReg_7),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~45_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~45 .extended_lut = "off";
defparam \sr~45 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~45 .shared_arith = "off";

cyclonev_lcell_comb \sr~46 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!sr_17),
	.datad(!MonDReg_15),
	.datae(!break_readreg_15),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~46_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~46 .extended_lut = "off";
defparam \sr~46 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~46 .shared_arith = "off";

cyclonev_lcell_comb \sr~47 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!MonDReg_8),
	.datad(!sr_10),
	.datae(!break_readreg_8),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~47_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~47 .extended_lut = "off";
defparam \sr~47 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~47 .shared_arith = "off";

cyclonev_lcell_comb \sr~48 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!MonDReg_9),
	.datad(!sr_11),
	.datae(!break_readreg_9),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~48_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~48 .extended_lut = "off";
defparam \sr~48 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~48 .shared_arith = "off";

cyclonev_lcell_comb \sr~49 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!MonDReg_10),
	.datad(!sr_12),
	.datae(!break_readreg_10),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~49_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~49 .extended_lut = "off";
defparam \sr~49 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~49 .shared_arith = "off";

cyclonev_lcell_comb \sr~52 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!MonDReg_12),
	.datad(!sr_14),
	.datae(!break_readreg_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~52_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~52 .extended_lut = "off";
defparam \sr~52 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~52 .shared_arith = "off";

cyclonev_lcell_comb \sr~53 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!MonDReg_13),
	.datad(!sr_15),
	.datae(!break_readreg_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~53_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~53 .extended_lut = "off";
defparam \sr~53 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~53 .shared_arith = "off";

cyclonev_lcell_comb \sr~54 (
	.dataa(!virtual_state_sdr),
	.datab(!irf_reg_1_1),
	.datac(!MonDReg_11),
	.datad(!sr_13),
	.datae(!break_readreg_11),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~54_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~54 .extended_lut = "off";
defparam \sr~54 .lut_mask = 64'h6FFFFFFF6FFFFFFF;
defparam \sr~54 .shared_arith = "off";

cyclonev_lcell_comb \sr~5 (
	.dataa(!sr_0),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!state_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~5 .extended_lut = "off";
defparam \sr~5 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \sr~5 .shared_arith = "off";

cyclonev_lcell_comb \sr~6 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!state_3),
	.datad(!\the_altera_std_synchronizer2|dreg[0]~q ),
	.datae(!irf_reg_0_1),
	.dataf(!irf_reg_1_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~6 .extended_lut = "off";
defparam \sr~6 .lut_mask = 64'hFFFFFFFFFFFFBFFF;
defparam \sr~6 .shared_arith = "off";

dffeas \DRsize.000 (
	.clk(altera_internal_jtag),
	.d(vcc),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.000~q ),
	.prn(vcc));
defparam \DRsize.000 .is_wysiwyg = "true";
defparam \DRsize.000 .power_up = "low";

cyclonev_lcell_comb \sr~7 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr~5_combout ),
	.datac(!\sr~6_combout ),
	.datad(!sr_1),
	.datae(!\DRsize.000~q ),
	.dataf(!altera_internal_jtag1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~7 .extended_lut = "off";
defparam \sr~7 .lut_mask = 64'h7FFFBFFFFFFFFFFF;
defparam \sr~7 .shared_arith = "off";

cyclonev_lcell_comb \sr~14 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!sr_37),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~14 .extended_lut = "off";
defparam \sr~14 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~14 .shared_arith = "off";

cyclonev_lcell_comb \sr[36]~15 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!state_3),
	.datae(!irf_reg_0_1),
	.dataf(!irf_reg_1_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[36]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[36]~15 .extended_lut = "off";
defparam \sr[36]~15 .lut_mask = 64'hDFFFFFFFFFFFDFFF;
defparam \sr[36]~15 .shared_arith = "off";

cyclonev_lcell_comb \sr~16 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(!altera_internal_jtag1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~16 .extended_lut = "off";
defparam \sr~16 .lut_mask = 64'hDFFFDFFFDFFFDFFF;
defparam \sr~16 .shared_arith = "off";

cyclonev_lcell_comb \Mux37~0 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_1_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Mux37~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Mux37~0 .extended_lut = "off";
defparam \Mux37~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \Mux37~0 .shared_arith = "off";

dffeas \DRsize.100 (
	.clk(altera_internal_jtag),
	.d(\Mux37~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.100~q ),
	.prn(vcc));
defparam \DRsize.100 .is_wysiwyg = "true";
defparam \DRsize.100 .power_up = "low";

cyclonev_lcell_comb \sr~56 (
	.dataa(!virtual_state_cdr),
	.datab(!sr_35),
	.datac(!irf_reg_0_1),
	.datad(!irf_reg_1_1),
	.datae(!\the_altera_std_synchronizer1|dreg[0]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~56_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~56 .extended_lut = "off";
defparam \sr~56 .lut_mask = 64'hB77BFFFFB77BFFFF;
defparam \sr~56 .shared_arith = "off";

cyclonev_lcell_comb \sr~17 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_36),
	.datad(!\DRsize.100~q ),
	.datae(!\sr~56_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~17 .extended_lut = "off";
defparam \sr~17 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~17 .shared_arith = "off";

cyclonev_lcell_comb \sr~18 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_35),
	.datad(!monitor_error),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~18 .extended_lut = "off";
defparam \sr~18 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~18 .shared_arith = "off";

cyclonev_lcell_comb \sr[23]~32 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!state_3),
	.datad(!irf_reg_0_1),
	.datae(!irf_reg_1_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[23]~32_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[23]~32 .extended_lut = "off";
defparam \sr[23]~32 .lut_mask = 64'hFFFFFFBFFFFFFFBF;
defparam \sr[23]~32 .shared_arith = "off";

cyclonev_lcell_comb \sr~33 (
	.dataa(!irf_reg_1_1),
	.datab(!MonDReg_30),
	.datac(!break_readreg_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~33_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~33 .extended_lut = "off";
defparam \sr~33 .lut_mask = 64'h2727272727272727;
defparam \sr~33 .shared_arith = "off";

cyclonev_lcell_comb \sr~34 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!state_3),
	.datad(!irf_reg_0_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~34_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~34 .extended_lut = "off";
defparam \sr~34 .lut_mask = 64'hFFBFFFBFFFBFFFBF;
defparam \sr~34 .shared_arith = "off";

cyclonev_lcell_comb \sr~35 (
	.dataa(!virtual_state_sdr),
	.datab(!\sr[23]~32_combout ),
	.datac(!sr_31),
	.datad(!sr_32),
	.datae(!\sr~33_combout ),
	.dataf(!\sr~34_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~35_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~35 .extended_lut = "off";
defparam \sr~35 .lut_mask = 64'h8DFFFFFFFFFFFFFF;
defparam \sr~35 .shared_arith = "off";

cyclonev_lcell_comb \sr~37 (
	.dataa(!virtual_state_sdr),
	.datab(!\Mux37~0_combout ),
	.datac(!sr_34),
	.datad(!resetlatch),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~37_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~37 .extended_lut = "off";
defparam \sr~37 .lut_mask = 64'h27FF27FF27FF27FF;
defparam \sr~37 .shared_arith = "off";

cyclonev_lcell_comb \sr~41 (
	.dataa(!irf_reg_1_1),
	.datab(!break_readreg_6),
	.datac(!MonDReg_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~41_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~41 .extended_lut = "off";
defparam \sr~41 .lut_mask = 64'h2727272727272727;
defparam \sr~41 .shared_arith = "off";

cyclonev_lcell_comb \sr~42 (
	.dataa(!virtual_state_sdr),
	.datab(!virtual_state_cdr),
	.datac(!irf_reg_0_1),
	.datad(!sr_7),
	.datae(!sr_8),
	.dataf(!\sr~41_combout ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~42_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~42 .extended_lut = "off";
defparam \sr~42 .lut_mask = 64'hF6FFFFFFFFFFFFFF;
defparam \sr~42 .shared_arith = "off";

cyclonev_lcell_comb \sr[23]~55 (
	.dataa(!irf_reg_0_1),
	.datab(!irf_reg_1_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr[23]~55_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr[23]~55 .extended_lut = "off";
defparam \sr[23]~55 .lut_mask = 64'h7777777777777777;
defparam \sr[23]~55 .shared_arith = "off";

dffeas \DRsize.010 (
	.clk(altera_internal_jtag),
	.d(\sr[23]~55_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(virtual_state_uir),
	.q(\DRsize.010~q ),
	.prn(vcc));
defparam \DRsize.010 .is_wysiwyg = "true";
defparam \DRsize.010 .power_up = "low";

cyclonev_lcell_comb \sr~50 (
	.dataa(!virtual_state_cdr),
	.datab(!irf_reg_0_1),
	.datac(!irf_reg_1_1),
	.datad(!MonDReg_14),
	.datae(!sr_15),
	.dataf(!break_readreg_14),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~50_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~50 .extended_lut = "off";
defparam \sr~50 .lut_mask = 64'hDEFFFFFFFFFFFFFF;
defparam \sr~50 .shared_arith = "off";

cyclonev_lcell_comb \sr~51 (
	.dataa(!virtual_state_sdr),
	.datab(!altera_internal_jtag1),
	.datac(!sr_16),
	.datad(!\DRsize.010~q ),
	.datae(!\sr~50_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sr~51_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sr~51 .extended_lut = "off";
defparam \sr~51 .lut_mask = 64'h7FBFFFFF7FBFFFFF;
defparam \sr~51 .shared_arith = "off";

endmodule

module embedded_system_altera_std_synchronizer_2 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module embedded_system_altera_std_synchronizer_3 (
	dreg_0,
	din,
	clk)/* synthesis synthesis_greybox=1 */;
output 	dreg_0;
input 	din;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module embedded_system_sld_virtual_jtag_basic_1 (
	virtual_state_sdr,
	virtual_state_uir1,
	virtual_state_cdr1,
	virtual_state_udr,
	state_4,
	splitter_nodes_receive_0_3,
	virtual_ir_scan_reg,
	state_3,
	state_8)/* synthesis synthesis_greybox=1 */;
output 	virtual_state_sdr;
output 	virtual_state_uir1;
output 	virtual_state_cdr1;
output 	virtual_state_udr;
input 	state_4;
input 	splitter_nodes_receive_0_3;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cyclonev_lcell_comb \virtual_state_sdr~0 (
	.dataa(!state_4),
	.datab(!virtual_ir_scan_reg),
	.datac(!splitter_nodes_receive_0_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_sdr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_sdr~0 .extended_lut = "off";
defparam \virtual_state_sdr~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \virtual_state_sdr~0 .shared_arith = "off";

cyclonev_lcell_comb virtual_state_uir(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_uir1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_uir.extended_lut = "off";
defparam virtual_state_uir.lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam virtual_state_uir.shared_arith = "off";

cyclonev_lcell_comb virtual_state_cdr(
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!state_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_cdr1),
	.sumout(),
	.cout(),
	.shareout());
defparam virtual_state_cdr.extended_lut = "off";
defparam virtual_state_cdr.lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam virtual_state_cdr.shared_arith = "off";

cyclonev_lcell_comb \virtual_state_udr~0 (
	.dataa(!virtual_ir_scan_reg),
	.datab(!splitter_nodes_receive_0_3),
	.datac(!state_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(virtual_state_udr),
	.sumout(),
	.cout(),
	.shareout());
defparam \virtual_state_udr~0 .extended_lut = "off";
defparam \virtual_state_udr~0 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \virtual_state_udr~0 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_nios2_avalon_reg (
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	write,
	address_8,
	address_0,
	address_4,
	address_3,
	address_2,
	address_1,
	address_7,
	address_6,
	address_5,
	Equal0,
	debugaccess,
	take_action_ocireg,
	oci_single_step_mode1,
	writedata_3,
	oci_reg_readdata,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
input 	write;
input 	address_8;
input 	address_0;
input 	address_4;
input 	address_3;
input 	address_2;
input 	address_1;
input 	address_7;
input 	address_6;
input 	address_5;
output 	Equal0;
input 	debugaccess;
output 	take_action_ocireg;
output 	oci_single_step_mode1;
input 	writedata_3;
output 	oci_reg_readdata;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Equal0~0_combout ;
wire \Equal0~1_combout ;
wire \oci_single_step_mode~0_combout ;
wire \oci_ienable[17]~0_combout ;
wire \oci_ienable[17]~q ;


cyclonev_lcell_comb \Equal0~2 (
	.dataa(!address_0),
	.datab(!\Equal0~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(Equal0),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~2 .extended_lut = "off";
defparam \Equal0~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \Equal0~2 .shared_arith = "off";

cyclonev_lcell_comb \take_action_ocireg~0 (
	.dataa(!write),
	.datab(!Equal0),
	.datac(!debugaccess),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(take_action_ocireg),
	.sumout(),
	.cout(),
	.shareout());
defparam \take_action_ocireg~0 .extended_lut = "off";
defparam \take_action_ocireg~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \take_action_ocireg~0 .shared_arith = "off";

dffeas oci_single_step_mode(
	.clk(clk_clk),
	.d(\oci_single_step_mode~0_combout ),
	.asdata(vcc),
	.clrn(!hq3myc14108phmpo7y7qmhbp98hy0vq),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(oci_single_step_mode1),
	.prn(vcc));
defparam oci_single_step_mode.is_wysiwyg = "true";
defparam oci_single_step_mode.power_up = "low";

cyclonev_lcell_comb \oci_reg_readdata~0 (
	.dataa(!address_0),
	.datab(!\Equal0~1_combout ),
	.datac(!\oci_ienable[17]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(oci_reg_readdata),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_reg_readdata~0 .extended_lut = "off";
defparam \oci_reg_readdata~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \oci_reg_readdata~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~0 (
	.dataa(!address_8),
	.datab(!address_7),
	.datac(!address_6),
	.datad(!address_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~0 .extended_lut = "off";
defparam \Equal0~0 .lut_mask = 64'hFFFDFFFDFFFDFFFD;
defparam \Equal0~0 .shared_arith = "off";

cyclonev_lcell_comb \Equal0~1 (
	.dataa(!address_4),
	.datab(!address_3),
	.datac(!address_2),
	.datad(!address_1),
	.datae(!\Equal0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Equal0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Equal0~1 .extended_lut = "off";
defparam \Equal0~1 .lut_mask = 64'hFFFEFFFFFFFEFFFF;
defparam \Equal0~1 .shared_arith = "off";

cyclonev_lcell_comb \oci_single_step_mode~0 (
	.dataa(!take_action_ocireg),
	.datab(!oci_single_step_mode1),
	.datac(!writedata_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_single_step_mode~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_single_step_mode~0 .extended_lut = "off";
defparam \oci_single_step_mode~0 .lut_mask = 64'h2727272727272727;
defparam \oci_single_step_mode~0 .shared_arith = "off";

cyclonev_lcell_comb \oci_ienable[17]~0 (
	.dataa(!write),
	.datab(!address_0),
	.datac(!\Equal0~1_combout ),
	.datad(!debugaccess),
	.datae(!\oci_ienable[17]~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\oci_ienable[17]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \oci_ienable[17]~0 .extended_lut = "off";
defparam \oci_ienable[17]~0 .lut_mask = 64'h7FFFFFFF7FFFFFFF;
defparam \oci_ienable[17]~0 .shared_arith = "off";

dffeas \oci_ienable[17] (
	.clk(clk_clk),
	.d(\oci_ienable[17]~0_combout ),
	.asdata(vcc),
	.clrn(!hq3myc14108phmpo7y7qmhbp98hy0vq),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\oci_ienable[17]~q ),
	.prn(vcc));
defparam \oci_ienable[17] .is_wysiwyg = "true";
defparam \oci_ienable[17] .power_up = "low";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_nios2_oci_break (
	break_readreg_0,
	break_readreg_1,
	break_readreg_2,
	break_readreg_3,
	break_readreg_24,
	break_readreg_4,
	break_readreg_20,
	break_readreg_19,
	break_readreg_16,
	break_readreg_25,
	break_readreg_5,
	break_readreg_26,
	break_readreg_27,
	break_readreg_28,
	break_readreg_29,
	break_readreg_30,
	break_readreg_31,
	break_readreg_21,
	break_readreg_18,
	break_readreg_17,
	break_readreg_6,
	break_readreg_22,
	break_readreg_23,
	break_readreg_7,
	break_readreg_15,
	break_readreg_8,
	break_readreg_9,
	break_readreg_10,
	break_readreg_14,
	break_readreg_12,
	break_readreg_13,
	break_readreg_11,
	jdo_0,
	jdo_36,
	jdo_37,
	ir_1,
	ir_0,
	enable_action_strobe,
	jdo_3,
	jdo_25,
	jdo_1,
	jdo_4,
	jdo_21,
	jdo_20,
	jdo_17,
	jdo_2,
	jdo_5,
	jdo_27,
	jdo_26,
	jdo_28,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_19,
	jdo_18,
	jdo_6,
	jdo_24,
	jdo_7,
	jdo_23,
	jdo_22,
	jdo_16,
	jdo_8,
	jdo_9,
	jdo_10,
	jdo_15,
	jdo_13,
	jdo_14,
	jdo_12,
	jdo_11,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	break_readreg_0;
output 	break_readreg_1;
output 	break_readreg_2;
output 	break_readreg_3;
output 	break_readreg_24;
output 	break_readreg_4;
output 	break_readreg_20;
output 	break_readreg_19;
output 	break_readreg_16;
output 	break_readreg_25;
output 	break_readreg_5;
output 	break_readreg_26;
output 	break_readreg_27;
output 	break_readreg_28;
output 	break_readreg_29;
output 	break_readreg_30;
output 	break_readreg_31;
output 	break_readreg_21;
output 	break_readreg_18;
output 	break_readreg_17;
output 	break_readreg_6;
output 	break_readreg_22;
output 	break_readreg_23;
output 	break_readreg_7;
output 	break_readreg_15;
output 	break_readreg_8;
output 	break_readreg_9;
output 	break_readreg_10;
output 	break_readreg_14;
output 	break_readreg_12;
output 	break_readreg_13;
output 	break_readreg_11;
input 	jdo_0;
input 	jdo_36;
input 	jdo_37;
input 	ir_1;
input 	ir_0;
input 	enable_action_strobe;
input 	jdo_3;
input 	jdo_25;
input 	jdo_1;
input 	jdo_4;
input 	jdo_21;
input 	jdo_20;
input 	jdo_17;
input 	jdo_2;
input 	jdo_5;
input 	jdo_27;
input 	jdo_26;
input 	jdo_28;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_19;
input 	jdo_18;
input 	jdo_6;
input 	jdo_24;
input 	jdo_7;
input 	jdo_23;
input 	jdo_22;
input 	jdo_16;
input 	jdo_8;
input 	jdo_9;
input 	jdo_10;
input 	jdo_15;
input 	jdo_13;
input 	jdo_14;
input 	jdo_12;
input 	jdo_11;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \break_readreg[4]~0_combout ;
wire \break_readreg[4]~1_combout ;


dffeas \break_readreg[0] (
	.clk(clk_clk),
	.d(jdo_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_0),
	.prn(vcc));
defparam \break_readreg[0] .is_wysiwyg = "true";
defparam \break_readreg[0] .power_up = "low";

dffeas \break_readreg[1] (
	.clk(clk_clk),
	.d(jdo_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_1),
	.prn(vcc));
defparam \break_readreg[1] .is_wysiwyg = "true";
defparam \break_readreg[1] .power_up = "low";

dffeas \break_readreg[2] (
	.clk(clk_clk),
	.d(jdo_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_2),
	.prn(vcc));
defparam \break_readreg[2] .is_wysiwyg = "true";
defparam \break_readreg[2] .power_up = "low";

dffeas \break_readreg[3] (
	.clk(clk_clk),
	.d(jdo_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_3),
	.prn(vcc));
defparam \break_readreg[3] .is_wysiwyg = "true";
defparam \break_readreg[3] .power_up = "low";

dffeas \break_readreg[24] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_24),
	.prn(vcc));
defparam \break_readreg[24] .is_wysiwyg = "true";
defparam \break_readreg[24] .power_up = "low";

dffeas \break_readreg[4] (
	.clk(clk_clk),
	.d(jdo_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_4),
	.prn(vcc));
defparam \break_readreg[4] .is_wysiwyg = "true";
defparam \break_readreg[4] .power_up = "low";

dffeas \break_readreg[20] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_20),
	.prn(vcc));
defparam \break_readreg[20] .is_wysiwyg = "true";
defparam \break_readreg[20] .power_up = "low";

dffeas \break_readreg[19] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_19),
	.prn(vcc));
defparam \break_readreg[19] .is_wysiwyg = "true";
defparam \break_readreg[19] .power_up = "low";

dffeas \break_readreg[16] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_16),
	.prn(vcc));
defparam \break_readreg[16] .is_wysiwyg = "true";
defparam \break_readreg[16] .power_up = "low";

dffeas \break_readreg[25] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_25),
	.prn(vcc));
defparam \break_readreg[25] .is_wysiwyg = "true";
defparam \break_readreg[25] .power_up = "low";

dffeas \break_readreg[5] (
	.clk(clk_clk),
	.d(jdo_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_5),
	.prn(vcc));
defparam \break_readreg[5] .is_wysiwyg = "true";
defparam \break_readreg[5] .power_up = "low";

dffeas \break_readreg[26] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_26),
	.prn(vcc));
defparam \break_readreg[26] .is_wysiwyg = "true";
defparam \break_readreg[26] .power_up = "low";

dffeas \break_readreg[27] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_27),
	.prn(vcc));
defparam \break_readreg[27] .is_wysiwyg = "true";
defparam \break_readreg[27] .power_up = "low";

dffeas \break_readreg[28] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_28),
	.prn(vcc));
defparam \break_readreg[28] .is_wysiwyg = "true";
defparam \break_readreg[28] .power_up = "low";

dffeas \break_readreg[29] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_29),
	.prn(vcc));
defparam \break_readreg[29] .is_wysiwyg = "true";
defparam \break_readreg[29] .power_up = "low";

dffeas \break_readreg[30] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_30),
	.prn(vcc));
defparam \break_readreg[30] .is_wysiwyg = "true";
defparam \break_readreg[30] .power_up = "low";

dffeas \break_readreg[31] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_31),
	.prn(vcc));
defparam \break_readreg[31] .is_wysiwyg = "true";
defparam \break_readreg[31] .power_up = "low";

dffeas \break_readreg[21] (
	.clk(clk_clk),
	.d(jdo_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_21),
	.prn(vcc));
defparam \break_readreg[21] .is_wysiwyg = "true";
defparam \break_readreg[21] .power_up = "low";

dffeas \break_readreg[18] (
	.clk(clk_clk),
	.d(jdo_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_18),
	.prn(vcc));
defparam \break_readreg[18] .is_wysiwyg = "true";
defparam \break_readreg[18] .power_up = "low";

dffeas \break_readreg[17] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_17),
	.prn(vcc));
defparam \break_readreg[17] .is_wysiwyg = "true";
defparam \break_readreg[17] .power_up = "low";

dffeas \break_readreg[6] (
	.clk(clk_clk),
	.d(jdo_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_6),
	.prn(vcc));
defparam \break_readreg[6] .is_wysiwyg = "true";
defparam \break_readreg[6] .power_up = "low";

dffeas \break_readreg[22] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_22),
	.prn(vcc));
defparam \break_readreg[22] .is_wysiwyg = "true";
defparam \break_readreg[22] .power_up = "low";

dffeas \break_readreg[23] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_23),
	.prn(vcc));
defparam \break_readreg[23] .is_wysiwyg = "true";
defparam \break_readreg[23] .power_up = "low";

dffeas \break_readreg[7] (
	.clk(clk_clk),
	.d(jdo_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_7),
	.prn(vcc));
defparam \break_readreg[7] .is_wysiwyg = "true";
defparam \break_readreg[7] .power_up = "low";

dffeas \break_readreg[15] (
	.clk(clk_clk),
	.d(jdo_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_15),
	.prn(vcc));
defparam \break_readreg[15] .is_wysiwyg = "true";
defparam \break_readreg[15] .power_up = "low";

dffeas \break_readreg[8] (
	.clk(clk_clk),
	.d(jdo_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_8),
	.prn(vcc));
defparam \break_readreg[8] .is_wysiwyg = "true";
defparam \break_readreg[8] .power_up = "low";

dffeas \break_readreg[9] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_9),
	.prn(vcc));
defparam \break_readreg[9] .is_wysiwyg = "true";
defparam \break_readreg[9] .power_up = "low";

dffeas \break_readreg[10] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_10),
	.prn(vcc));
defparam \break_readreg[10] .is_wysiwyg = "true";
defparam \break_readreg[10] .power_up = "low";

dffeas \break_readreg[14] (
	.clk(clk_clk),
	.d(jdo_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_14),
	.prn(vcc));
defparam \break_readreg[14] .is_wysiwyg = "true";
defparam \break_readreg[14] .power_up = "low";

dffeas \break_readreg[12] (
	.clk(clk_clk),
	.d(jdo_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_12),
	.prn(vcc));
defparam \break_readreg[12] .is_wysiwyg = "true";
defparam \break_readreg[12] .power_up = "low";

dffeas \break_readreg[13] (
	.clk(clk_clk),
	.d(jdo_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_13),
	.prn(vcc));
defparam \break_readreg[13] .is_wysiwyg = "true";
defparam \break_readreg[13] .power_up = "low";

dffeas \break_readreg[11] (
	.clk(clk_clk),
	.d(jdo_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\break_readreg[4]~1_combout ),
	.sload(gnd),
	.ena(\break_readreg[4]~0_combout ),
	.q(break_readreg_11),
	.prn(vcc));
defparam \break_readreg[11] .is_wysiwyg = "true";
defparam \break_readreg[11] .power_up = "low";

cyclonev_lcell_comb \break_readreg[4]~0 (
	.dataa(!ir_1),
	.datab(!ir_0),
	.datac(!enable_action_strobe),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[4]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[4]~0 .extended_lut = "off";
defparam \break_readreg[4]~0 .lut_mask = 64'hDFDFDFDFDFDFDFDF;
defparam \break_readreg[4]~0 .shared_arith = "off";

cyclonev_lcell_comb \break_readreg[4]~1 (
	.dataa(!jdo_36),
	.datab(!jdo_37),
	.datac(!\break_readreg[4]~0_combout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_readreg[4]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_readreg[4]~1 .extended_lut = "off";
defparam \break_readreg[4]~1 .lut_mask = 64'hEFEFEFEFEFEFEFEF;
defparam \break_readreg[4]~1 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_nios2_oci_debug (
	hq3myc14108phmpo7y7qmhbp98hy0vq,
	monitor_ready1,
	jtag_break1,
	take_action_ocimem_a,
	jdo_34,
	take_action_ocimem_a1,
	jdo_25,
	writedata_0,
	take_action_ocireg,
	jdo_21,
	jdo_20,
	writedata_1,
	jdo_19,
	jdo_18,
	monitor_error1,
	resetrequest1,
	jdo_24,
	resetlatch1,
	jdo_23,
	jdo_22,
	monitor_go1,
	state_1,
	clk_clk)/* synthesis synthesis_greybox=1 */;
input 	hq3myc14108phmpo7y7qmhbp98hy0vq;
output 	monitor_ready1;
output 	jtag_break1;
input 	take_action_ocimem_a;
input 	jdo_34;
input 	take_action_ocimem_a1;
input 	jdo_25;
input 	writedata_0;
input 	take_action_ocireg;
input 	jdo_21;
input 	jdo_20;
input 	writedata_1;
input 	jdo_19;
input 	jdo_18;
output 	monitor_error1;
output 	resetrequest1;
input 	jdo_24;
output 	resetlatch1;
input 	jdo_23;
input 	jdo_22;
output 	monitor_go1;
input 	state_1;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \the_altera_std_synchronizer|dreg[0]~q ;
wire \monitor_ready~0_combout ;
wire \break_on_reset~0_combout ;
wire \break_on_reset~q ;
wire \jtag_break~0_combout ;
wire \monitor_error~0_combout ;
wire \resetlatch~0_combout ;
wire \monitor_go~0_combout ;


embedded_system_altera_std_synchronizer_4 the_altera_std_synchronizer(
	.din(hq3myc14108phmpo7y7qmhbp98hy0vq),
	.dreg_0(\the_altera_std_synchronizer|dreg[0]~q ),
	.clk(clk_clk));

dffeas monitor_ready(
	.clk(clk_clk),
	.d(\monitor_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_ready1),
	.prn(vcc));
defparam monitor_ready.is_wysiwyg = "true";
defparam monitor_ready.power_up = "low";

dffeas jtag_break(
	.clk(clk_clk),
	.d(\jtag_break~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(jtag_break1),
	.prn(vcc));
defparam jtag_break.is_wysiwyg = "true";
defparam jtag_break.power_up = "low";

dffeas monitor_error(
	.clk(clk_clk),
	.d(\monitor_error~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_error1),
	.prn(vcc));
defparam monitor_error.is_wysiwyg = "true";
defparam monitor_error.power_up = "low";

dffeas resetrequest(
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a1),
	.q(resetrequest1),
	.prn(vcc));
defparam resetrequest.is_wysiwyg = "true";
defparam resetrequest.power_up = "low";

dffeas resetlatch(
	.clk(clk_clk),
	.d(\resetlatch~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(resetlatch1),
	.prn(vcc));
defparam resetlatch.is_wysiwyg = "true";
defparam resetlatch.power_up = "low";

dffeas monitor_go(
	.clk(clk_clk),
	.d(\monitor_go~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(monitor_go1),
	.prn(vcc));
defparam monitor_go.is_wysiwyg = "true";
defparam monitor_go.power_up = "low";

cyclonev_lcell_comb \monitor_ready~0 (
	.dataa(!monitor_ready1),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_25),
	.datad(!writedata_0),
	.datae(!take_action_ocireg),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_ready~0 .extended_lut = "off";
defparam \monitor_ready~0 .lut_mask = 64'hFDFFFFFFFDFFFFFF;
defparam \monitor_ready~0 .shared_arith = "off";

cyclonev_lcell_comb \break_on_reset~0 (
	.dataa(!\break_on_reset~q ),
	.datab(!jdo_19),
	.datac(!jdo_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\break_on_reset~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \break_on_reset~0 .extended_lut = "off";
defparam \break_on_reset~0 .lut_mask = 64'hF7F7F7F7F7F7F7F7;
defparam \break_on_reset~0 .shared_arith = "off";

dffeas break_on_reset(
	.clk(clk_clk),
	.d(\break_on_reset~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(take_action_ocimem_a1),
	.q(\break_on_reset~q ),
	.prn(vcc));
defparam break_on_reset.is_wysiwyg = "true";
defparam break_on_reset.power_up = "low";

cyclonev_lcell_comb \jtag_break~0 (
	.dataa(!jtag_break1),
	.datab(!take_action_ocimem_a1),
	.datac(!jdo_21),
	.datad(!jdo_20),
	.datae(!\break_on_reset~q ),
	.dataf(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_break~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_break~0 .extended_lut = "off";
defparam \jtag_break~0 .lut_mask = 64'hFF7FFFFFFFDFFFFF;
defparam \jtag_break~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_error~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!jdo_25),
	.datac(!take_action_ocireg),
	.datad(!writedata_1),
	.datae(!monitor_error1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_error~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_error~0 .extended_lut = "off";
defparam \monitor_error~0 .lut_mask = 64'hEFFFFFFFEFFFFFFF;
defparam \monitor_error~0 .shared_arith = "off";

cyclonev_lcell_comb \resetlatch~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!\the_altera_std_synchronizer|dreg[0]~q ),
	.datac(!jdo_24),
	.datad(!resetlatch1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\resetlatch~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \resetlatch~0 .extended_lut = "off";
defparam \resetlatch~0 .lut_mask = 64'hFBFFFBFFFBFFFBFF;
defparam \resetlatch~0 .shared_arith = "off";

cyclonev_lcell_comb \monitor_go~0 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_34),
	.datac(!jdo_23),
	.datad(!monitor_go1),
	.datae(!state_1),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\monitor_go~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \monitor_go~0 .extended_lut = "off";
defparam \monitor_go~0 .lut_mask = 64'hFFFF7FFFFFFF7FFF;
defparam \monitor_go~0 .shared_arith = "off";

endmodule

module embedded_system_altera_std_synchronizer_4 (
	din,
	dreg_0,
	clk)/* synthesis synthesis_greybox=1 */;
input 	din;
output 	dreg_0;
input 	clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \din_s1~q ;


dffeas \dreg[0] (
	.clk(clk),
	.d(\din_s1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(dreg_0),
	.prn(vcc));
defparam \dreg[0] .is_wysiwyg = "true";
defparam \dreg[0] .power_up = "low";

dffeas din_s1(
	.clk(clk),
	.d(din),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\din_s1~q ),
	.prn(vcc));
defparam din_s1.is_wysiwyg = "true";
defparam din_s1.power_up = "low";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_nios2_ocimem (
	MonDReg_0,
	q_a_0,
	q_a_1,
	q_a_2,
	MonDReg_24,
	MonDReg_4,
	q_a_3,
	MonDReg_20,
	MonDReg_19,
	MonDReg_16,
	MonDReg_25,
	q_a_24,
	q_a_4,
	MonDReg_26,
	MonDReg_27,
	MonDReg_28,
	MonDReg_30,
	MonDReg_31,
	MonDReg_21,
	q_a_20,
	q_a_19,
	MonDReg_17,
	q_a_16,
	q_a_25,
	MonDReg_6,
	q_a_5,
	q_a_26,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	MonDReg_22,
	q_a_21,
	q_a_18,
	q_a_17,
	q_a_10,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_13,
	q_a_12,
	q_a_11,
	q_a_9,
	q_a_8,
	q_a_6,
	q_a_14,
	q_a_22,
	MonDReg_23,
	MonDReg_7,
	MonDReg_15,
	MonDReg_13,
	MonDReg_14,
	waitrequest1,
	MonDReg_1,
	jdo_3,
	take_action_ocimem_a,
	jdo_35,
	take_action_ocimem_b,
	write,
	address_8,
	read,
	take_action_ocimem_a1,
	jdo_34,
	take_action_ocimem_a2,
	jdo_25,
	writedata_0,
	address_0,
	address_4,
	address_3,
	address_2,
	address_1,
	address_7,
	address_6,
	address_5,
	debugaccess,
	MonDReg_2,
	jdo_4,
	r_early_rst,
	byteenable_0,
	jdo_21,
	jdo_20,
	jdo_17,
	MonDReg_3,
	jdo_5,
	writedata_1,
	jdo_27,
	jdo_26,
	jdo_28,
	jdo_29,
	jdo_30,
	jdo_31,
	jdo_32,
	jdo_33,
	writedata_3,
	jdo_19,
	jdo_18,
	jdo_6,
	writedata_2,
	jdo_24,
	MonDReg_5,
	jdo_7,
	MonDReg_29,
	jdo_23,
	jdo_22,
	MonDReg_18,
	jdo_16,
	writedata_24,
	byteenable_3,
	jdo_8,
	writedata_4,
	writedata_20,
	byteenable_2,
	writedata_19,
	writedata_16,
	writedata_25,
	jdo_9,
	writedata_5,
	writedata_26,
	writedata_27,
	writedata_28,
	writedata_29,
	writedata_30,
	writedata_31,
	writedata_21,
	writedata_18,
	writedata_17,
	MonDReg_10,
	writedata_10,
	byteenable_1,
	writedata_7,
	writedata_23,
	writedata_15,
	writedata_13,
	MonDReg_12,
	writedata_12,
	MonDReg_11,
	writedata_11,
	MonDReg_9,
	writedata_9,
	MonDReg_8,
	writedata_8,
	writedata_6,
	writedata_14,
	writedata_22,
	jdo_10,
	jdo_15,
	jdo_13,
	jdo_14,
	jdo_12,
	jdo_11,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	MonDReg_0;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	MonDReg_24;
output 	MonDReg_4;
output 	q_a_3;
output 	MonDReg_20;
output 	MonDReg_19;
output 	MonDReg_16;
output 	MonDReg_25;
output 	q_a_24;
output 	q_a_4;
output 	MonDReg_26;
output 	MonDReg_27;
output 	MonDReg_28;
output 	MonDReg_30;
output 	MonDReg_31;
output 	MonDReg_21;
output 	q_a_20;
output 	q_a_19;
output 	MonDReg_17;
output 	q_a_16;
output 	q_a_25;
output 	MonDReg_6;
output 	q_a_5;
output 	q_a_26;
output 	q_a_27;
output 	q_a_28;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
output 	MonDReg_22;
output 	q_a_21;
output 	q_a_18;
output 	q_a_17;
output 	q_a_10;
output 	q_a_7;
output 	q_a_23;
output 	q_a_15;
output 	q_a_13;
output 	q_a_12;
output 	q_a_11;
output 	q_a_9;
output 	q_a_8;
output 	q_a_6;
output 	q_a_14;
output 	q_a_22;
output 	MonDReg_23;
output 	MonDReg_7;
output 	MonDReg_15;
output 	MonDReg_13;
output 	MonDReg_14;
output 	waitrequest1;
output 	MonDReg_1;
input 	jdo_3;
input 	take_action_ocimem_a;
input 	jdo_35;
input 	take_action_ocimem_b;
input 	write;
input 	address_8;
input 	read;
input 	take_action_ocimem_a1;
input 	jdo_34;
input 	take_action_ocimem_a2;
input 	jdo_25;
input 	writedata_0;
input 	address_0;
input 	address_4;
input 	address_3;
input 	address_2;
input 	address_1;
input 	address_7;
input 	address_6;
input 	address_5;
input 	debugaccess;
output 	MonDReg_2;
input 	jdo_4;
input 	r_early_rst;
input 	byteenable_0;
input 	jdo_21;
input 	jdo_20;
input 	jdo_17;
output 	MonDReg_3;
input 	jdo_5;
input 	writedata_1;
input 	jdo_27;
input 	jdo_26;
input 	jdo_28;
input 	jdo_29;
input 	jdo_30;
input 	jdo_31;
input 	jdo_32;
input 	jdo_33;
input 	writedata_3;
input 	jdo_19;
input 	jdo_18;
input 	jdo_6;
input 	writedata_2;
input 	jdo_24;
output 	MonDReg_5;
input 	jdo_7;
output 	MonDReg_29;
input 	jdo_23;
input 	jdo_22;
output 	MonDReg_18;
input 	jdo_16;
input 	writedata_24;
input 	byteenable_3;
input 	jdo_8;
input 	writedata_4;
input 	writedata_20;
input 	byteenable_2;
input 	writedata_19;
input 	writedata_16;
input 	writedata_25;
input 	jdo_9;
input 	writedata_5;
input 	writedata_26;
input 	writedata_27;
input 	writedata_28;
input 	writedata_29;
input 	writedata_30;
input 	writedata_31;
input 	writedata_21;
input 	writedata_18;
input 	writedata_17;
output 	MonDReg_10;
input 	writedata_10;
input 	byteenable_1;
input 	writedata_7;
input 	writedata_23;
input 	writedata_15;
input 	writedata_13;
output 	MonDReg_12;
input 	writedata_12;
output 	MonDReg_11;
input 	writedata_11;
output 	MonDReg_9;
input 	writedata_9;
output 	MonDReg_8;
input 	writedata_8;
input 	writedata_6;
input 	writedata_14;
input 	writedata_22;
input 	jdo_10;
input 	jdo_15;
input 	jdo_13;
input 	jdo_14;
input 	jdo_12;
input 	jdo_11;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \jtag_ram_wr~q ;
wire \ociram_wr_en~0_combout ;
wire \ociram_reset_req~combout ;
wire \ociram_wr_data[0]~0_combout ;
wire \ociram_addr[0]~0_combout ;
wire \ociram_addr[1]~1_combout ;
wire \ociram_addr[2]~2_combout ;
wire \ociram_addr[3]~3_combout ;
wire \ociram_addr[4]~4_combout ;
wire \ociram_addr[5]~5_combout ;
wire \ociram_addr[6]~6_combout ;
wire \ociram_addr[7]~7_combout ;
wire \ociram_byteenable[0]~0_combout ;
wire \ociram_wr_data[1]~1_combout ;
wire \jtag_ram_wr~0_combout ;
wire \ociram_wr_data[2]~2_combout ;
wire \ociram_wr_data[3]~3_combout ;
wire \ociram_wr_data[24]~4_combout ;
wire \ociram_byteenable[3]~1_combout ;
wire \ociram_wr_data[4]~5_combout ;
wire \ociram_wr_data[20]~6_combout ;
wire \ociram_byteenable[2]~2_combout ;
wire \ociram_wr_data[19]~7_combout ;
wire \ociram_wr_data[16]~8_combout ;
wire \ociram_wr_data[25]~9_combout ;
wire \ociram_wr_data[5]~10_combout ;
wire \ociram_wr_data[26]~11_combout ;
wire \ociram_wr_data[27]~12_combout ;
wire \ociram_wr_data[28]~13_combout ;
wire \ociram_wr_data[29]~14_combout ;
wire \ociram_wr_data[30]~15_combout ;
wire \ociram_wr_data[31]~16_combout ;
wire \ociram_wr_data[21]~17_combout ;
wire \ociram_wr_data[18]~18_combout ;
wire \ociram_wr_data[17]~19_combout ;
wire \ociram_wr_data[10]~20_combout ;
wire \ociram_byteenable[1]~3_combout ;
wire \ociram_wr_data[7]~21_combout ;
wire \ociram_wr_data[23]~22_combout ;
wire \ociram_wr_data[15]~23_combout ;
wire \ociram_wr_data[13]~24_combout ;
wire \ociram_wr_data[12]~25_combout ;
wire \ociram_wr_data[11]~26_combout ;
wire \ociram_wr_data[9]~27_combout ;
wire \ociram_wr_data[8]~28_combout ;
wire \ociram_wr_data[6]~29_combout ;
wire \ociram_wr_data[14]~30_combout ;
wire \ociram_wr_data[22]~31_combout ;
wire \Add0~1_wirecell_combout ;
wire \MonAReg[10]~q ;
wire \Add0~9_sumout ;
wire \MonAReg[2]~q ;
wire \Add0~10 ;
wire \Add0~5_sumout ;
wire \MonAReg[3]~q ;
wire \Add0~6 ;
wire \Add0~13_sumout ;
wire \MonAReg[4]~q ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \MonAReg[5]~q ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \MonAReg[6]~q ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \MonAReg[7]~q ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \MonAReg[8]~q ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \MonAReg[9]~q ;
wire \Add0~34 ;
wire \Add0~1_sumout ;
wire \jtag_ram_rd~0_combout ;
wire \jtag_ram_rd~q ;
wire \jtag_ram_rd_d1~q ;
wire \MonDReg[23]~0_combout ;
wire \jtag_rd~q ;
wire \jtag_rd_d1~q ;
wire \MonDReg[0]~1_combout ;
wire \jtag_ram_access~0_combout ;
wire \jtag_ram_access~q ;
wire \waitrequest~0_combout ;
wire \avalon_ociram_readdata_ready~0_combout ;
wire \avalon_ociram_readdata_ready~q ;
wire \waitrequest~1_combout ;
wire \MonDReg~2_combout ;
wire \MonDReg~3_combout ;
wire \MonDReg~4_combout ;
wire \MonDReg~5_combout ;
wire \MonDReg~6_combout ;
wire \MonDReg~27_combout ;
wire \MonDReg~23_combout ;
wire \MonDReg~19_combout ;
wire \MonDReg~7_combout ;
wire \MonDReg[12]~15_combout ;
wire \MonDReg[12]~8_combout ;
wire \MonDReg~9_combout ;
wire \MonDReg~10_combout ;
wire \MonDReg[8]~11_combout ;


embedded_system_embedded_system_nios2_qsys_0_ociram_sp_ram_module embedded_system_nios2_qsys_0_ociram_sp_ram(
	.q_a_0(q_a_0),
	.q_a_1(q_a_1),
	.q_a_2(q_a_2),
	.q_a_3(q_a_3),
	.q_a_24(q_a_24),
	.q_a_4(q_a_4),
	.q_a_20(q_a_20),
	.q_a_19(q_a_19),
	.q_a_16(q_a_16),
	.q_a_25(q_a_25),
	.q_a_5(q_a_5),
	.q_a_26(q_a_26),
	.q_a_27(q_a_27),
	.q_a_28(q_a_28),
	.q_a_29(q_a_29),
	.q_a_30(q_a_30),
	.q_a_31(q_a_31),
	.q_a_21(q_a_21),
	.q_a_18(q_a_18),
	.q_a_17(q_a_17),
	.q_a_10(q_a_10),
	.q_a_7(q_a_7),
	.q_a_23(q_a_23),
	.q_a_15(q_a_15),
	.q_a_13(q_a_13),
	.q_a_12(q_a_12),
	.q_a_11(q_a_11),
	.q_a_9(q_a_9),
	.q_a_8(q_a_8),
	.q_a_6(q_a_6),
	.q_a_14(q_a_14),
	.q_a_22(q_a_22),
	.ociram_wr_en(\ociram_wr_en~0_combout ),
	.ociram_reset_req(\ociram_reset_req~combout ),
	.ociram_wr_data_0(\ociram_wr_data[0]~0_combout ),
	.ociram_addr_0(\ociram_addr[0]~0_combout ),
	.ociram_addr_1(\ociram_addr[1]~1_combout ),
	.ociram_addr_2(\ociram_addr[2]~2_combout ),
	.ociram_addr_3(\ociram_addr[3]~3_combout ),
	.ociram_addr_4(\ociram_addr[4]~4_combout ),
	.ociram_addr_5(\ociram_addr[5]~5_combout ),
	.ociram_addr_6(\ociram_addr[6]~6_combout ),
	.ociram_addr_7(\ociram_addr[7]~7_combout ),
	.ociram_byteenable_0(\ociram_byteenable[0]~0_combout ),
	.ociram_wr_data_1(\ociram_wr_data[1]~1_combout ),
	.ociram_wr_data_2(\ociram_wr_data[2]~2_combout ),
	.ociram_wr_data_3(\ociram_wr_data[3]~3_combout ),
	.ociram_wr_data_24(\ociram_wr_data[24]~4_combout ),
	.ociram_byteenable_3(\ociram_byteenable[3]~1_combout ),
	.ociram_wr_data_4(\ociram_wr_data[4]~5_combout ),
	.ociram_wr_data_20(\ociram_wr_data[20]~6_combout ),
	.ociram_byteenable_2(\ociram_byteenable[2]~2_combout ),
	.ociram_wr_data_19(\ociram_wr_data[19]~7_combout ),
	.ociram_wr_data_16(\ociram_wr_data[16]~8_combout ),
	.ociram_wr_data_25(\ociram_wr_data[25]~9_combout ),
	.ociram_wr_data_5(\ociram_wr_data[5]~10_combout ),
	.ociram_wr_data_26(\ociram_wr_data[26]~11_combout ),
	.ociram_wr_data_27(\ociram_wr_data[27]~12_combout ),
	.ociram_wr_data_28(\ociram_wr_data[28]~13_combout ),
	.ociram_wr_data_29(\ociram_wr_data[29]~14_combout ),
	.ociram_wr_data_30(\ociram_wr_data[30]~15_combout ),
	.ociram_wr_data_31(\ociram_wr_data[31]~16_combout ),
	.ociram_wr_data_21(\ociram_wr_data[21]~17_combout ),
	.ociram_wr_data_18(\ociram_wr_data[18]~18_combout ),
	.ociram_wr_data_17(\ociram_wr_data[17]~19_combout ),
	.ociram_wr_data_10(\ociram_wr_data[10]~20_combout ),
	.ociram_byteenable_1(\ociram_byteenable[1]~3_combout ),
	.ociram_wr_data_7(\ociram_wr_data[7]~21_combout ),
	.ociram_wr_data_23(\ociram_wr_data[23]~22_combout ),
	.ociram_wr_data_15(\ociram_wr_data[15]~23_combout ),
	.ociram_wr_data_13(\ociram_wr_data[13]~24_combout ),
	.ociram_wr_data_12(\ociram_wr_data[12]~25_combout ),
	.ociram_wr_data_11(\ociram_wr_data[11]~26_combout ),
	.ociram_wr_data_9(\ociram_wr_data[9]~27_combout ),
	.ociram_wr_data_8(\ociram_wr_data[8]~28_combout ),
	.ociram_wr_data_6(\ociram_wr_data[6]~29_combout ),
	.ociram_wr_data_14(\ociram_wr_data[14]~30_combout ),
	.ociram_wr_data_22(\ociram_wr_data[22]~31_combout ),
	.clk_clk(clk_clk));

dffeas jtag_ram_wr(
	.clk(clk_clk),
	.d(\jtag_ram_wr~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_wr~q ),
	.prn(vcc));
defparam jtag_ram_wr.is_wysiwyg = "true";
defparam jtag_ram_wr.power_up = "low";

cyclonev_lcell_comb \ociram_wr_en~0 (
	.dataa(!write),
	.datab(!address_8),
	.datac(!\jtag_ram_access~q ),
	.datad(!debugaccess),
	.datae(!\jtag_ram_wr~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_en~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_en~0 .extended_lut = "off";
defparam \ociram_wr_en~0 .lut_mask = 64'hC5FFFFFFC5FFFFFF;
defparam \ociram_wr_en~0 .shared_arith = "off";

cyclonev_lcell_comb ociram_reset_req(
	.dataa(!\jtag_ram_access~q ),
	.datab(!r_early_rst),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_reset_req~combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam ociram_reset_req.extended_lut = "off";
defparam ociram_reset_req.lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam ociram_reset_req.shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[0]~0 (
	.dataa(!MonDReg_0),
	.datab(!\jtag_ram_access~q ),
	.datac(!writedata_0),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[0]~0 .extended_lut = "off";
defparam \ociram_wr_data[0]~0 .lut_mask = 64'h4747474747474747;
defparam \ociram_wr_data[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!address_0),
	.datac(!\MonAReg[2]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[0]~0 .extended_lut = "off";
defparam \ociram_addr[0]~0 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[1]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!address_1),
	.datac(!\MonAReg[3]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[1]~1 .extended_lut = "off";
defparam \ociram_addr[1]~1 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!address_2),
	.datac(!\MonAReg[4]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[2]~2 .extended_lut = "off";
defparam \ociram_addr[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[3]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!address_3),
	.datac(!\MonAReg[5]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[3]~3 .extended_lut = "off";
defparam \ociram_addr[3]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[4]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!address_4),
	.datac(!\MonAReg[6]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[4]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[4]~4 .extended_lut = "off";
defparam \ociram_addr[4]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[4]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[5]~5 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!address_5),
	.datac(!\MonAReg[7]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[5]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[5]~5 .extended_lut = "off";
defparam \ociram_addr[5]~5 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[5]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[6]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!address_6),
	.datac(!\MonAReg[8]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[6]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[6]~6 .extended_lut = "off";
defparam \ociram_addr[6]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[6]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_addr[7]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!address_7),
	.datac(!\MonAReg[9]~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_addr[7]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_addr[7]~7 .extended_lut = "off";
defparam \ociram_addr[7]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_addr[7]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[0]~0 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_0),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[0]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[0]~0 .extended_lut = "off";
defparam \ociram_byteenable[0]~0 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[0]~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[1]~1 (
	.dataa(!MonDReg_1),
	.datab(!\jtag_ram_access~q ),
	.datac(!writedata_1),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[1]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[1]~1 .extended_lut = "off";
defparam \ociram_wr_data[1]~1 .lut_mask = 64'h4747474747474747;
defparam \ociram_wr_data[1]~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_wr~0 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_35),
	.datac(!\jtag_ram_wr~q ),
	.datad(!\Add0~1_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_wr~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_wr~0 .extended_lut = "off";
defparam \jtag_ram_wr~0 .lut_mask = 64'h47FF47FF47FF47FF;
defparam \jtag_ram_wr~0 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_2),
	.datac(!writedata_2),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[2]~2 .extended_lut = "off";
defparam \ociram_wr_data[2]~2 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[3]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_3),
	.datac(!writedata_3),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[3]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[3]~3 .extended_lut = "off";
defparam \ociram_wr_data[3]~3 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[3]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[24]~4 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_24),
	.datac(!writedata_24),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[24]~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[24]~4 .extended_lut = "off";
defparam \ociram_wr_data[24]~4 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[24]~4 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[3]~1 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[3]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[3]~1 .extended_lut = "off";
defparam \ociram_byteenable[3]~1 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[3]~1 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[4]~5 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_4),
	.datac(!writedata_4),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[4]~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[4]~5 .extended_lut = "off";
defparam \ociram_wr_data[4]~5 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[4]~5 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[20]~6 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_20),
	.datac(!writedata_20),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[20]~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[20]~6 .extended_lut = "off";
defparam \ociram_wr_data[20]~6 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[20]~6 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[2]~2 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[2]~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[2]~2 .extended_lut = "off";
defparam \ociram_byteenable[2]~2 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[2]~2 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[19]~7 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_19),
	.datac(!writedata_19),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[19]~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[19]~7 .extended_lut = "off";
defparam \ociram_wr_data[19]~7 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[19]~7 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[16]~8 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_16),
	.datac(!writedata_16),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[16]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[16]~8 .extended_lut = "off";
defparam \ociram_wr_data[16]~8 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[16]~8 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[25]~9 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_25),
	.datac(!writedata_25),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[25]~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[25]~9 .extended_lut = "off";
defparam \ociram_wr_data[25]~9 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[25]~9 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[5]~10 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_5),
	.datac(!writedata_5),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[5]~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[5]~10 .extended_lut = "off";
defparam \ociram_wr_data[5]~10 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[5]~10 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[26]~11 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_26),
	.datac(!writedata_26),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[26]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[26]~11 .extended_lut = "off";
defparam \ociram_wr_data[26]~11 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[26]~11 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[27]~12 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_27),
	.datac(!writedata_27),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[27]~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[27]~12 .extended_lut = "off";
defparam \ociram_wr_data[27]~12 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[27]~12 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[28]~13 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_28),
	.datac(!writedata_28),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[28]~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[28]~13 .extended_lut = "off";
defparam \ociram_wr_data[28]~13 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[28]~13 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[29]~14 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_29),
	.datac(!writedata_29),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[29]~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[29]~14 .extended_lut = "off";
defparam \ociram_wr_data[29]~14 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[29]~14 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[30]~15 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_30),
	.datac(!writedata_30),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[30]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[30]~15 .extended_lut = "off";
defparam \ociram_wr_data[30]~15 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[30]~15 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[31]~16 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_31),
	.datac(!writedata_31),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[31]~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[31]~16 .extended_lut = "off";
defparam \ociram_wr_data[31]~16 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[31]~16 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[21]~17 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_21),
	.datac(!writedata_21),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[21]~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[21]~17 .extended_lut = "off";
defparam \ociram_wr_data[21]~17 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[21]~17 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[18]~18 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_18),
	.datac(!writedata_18),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[18]~18_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[18]~18 .extended_lut = "off";
defparam \ociram_wr_data[18]~18 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[18]~18 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[17]~19 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_17),
	.datac(!writedata_17),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[17]~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[17]~19 .extended_lut = "off";
defparam \ociram_wr_data[17]~19 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[17]~19 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[10]~20 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_10),
	.datac(!writedata_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[10]~20_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[10]~20 .extended_lut = "off";
defparam \ociram_wr_data[10]~20 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[10]~20 .shared_arith = "off";

cyclonev_lcell_comb \ociram_byteenable[1]~3 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!byteenable_1),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_byteenable[1]~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_byteenable[1]~3 .extended_lut = "off";
defparam \ociram_byteenable[1]~3 .lut_mask = 64'h7777777777777777;
defparam \ociram_byteenable[1]~3 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[7]~21 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_7),
	.datac(!writedata_7),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[7]~21_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[7]~21 .extended_lut = "off";
defparam \ociram_wr_data[7]~21 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[7]~21 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[23]~22 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_23),
	.datac(!writedata_23),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[23]~22_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[23]~22 .extended_lut = "off";
defparam \ociram_wr_data[23]~22 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[23]~22 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[15]~23 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_15),
	.datac(!writedata_15),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[15]~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[15]~23 .extended_lut = "off";
defparam \ociram_wr_data[15]~23 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[15]~23 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[13]~24 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_13),
	.datac(!writedata_13),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[13]~24_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[13]~24 .extended_lut = "off";
defparam \ociram_wr_data[13]~24 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[13]~24 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[12]~25 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_12),
	.datac(!writedata_12),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[12]~25_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[12]~25 .extended_lut = "off";
defparam \ociram_wr_data[12]~25 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[12]~25 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[11]~26 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_11),
	.datac(!writedata_11),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[11]~26_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[11]~26 .extended_lut = "off";
defparam \ociram_wr_data[11]~26 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[11]~26 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[9]~27 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_9),
	.datac(!writedata_9),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[9]~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[9]~27 .extended_lut = "off";
defparam \ociram_wr_data[9]~27 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[9]~27 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[8]~28 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_8),
	.datac(!writedata_8),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[8]~28_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[8]~28 .extended_lut = "off";
defparam \ociram_wr_data[8]~28 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[8]~28 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[6]~29 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_6),
	.datac(!writedata_6),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[6]~29_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[6]~29 .extended_lut = "off";
defparam \ociram_wr_data[6]~29 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[6]~29 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[14]~30 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_14),
	.datac(!writedata_14),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[14]~30_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[14]~30 .extended_lut = "off";
defparam \ociram_wr_data[14]~30 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[14]~30 .shared_arith = "off";

cyclonev_lcell_comb \ociram_wr_data[22]~31 (
	.dataa(!\jtag_ram_access~q ),
	.datab(!MonDReg_22),
	.datac(!writedata_22),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\ociram_wr_data[22]~31_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \ociram_wr_data[22]~31 .extended_lut = "off";
defparam \ociram_wr_data[22]~31 .lut_mask = 64'h2727272727272727;
defparam \ociram_wr_data[22]~31 .shared_arith = "off";

dffeas \MonDReg[0] (
	.clk(clk_clk),
	.d(jdo_3),
	.asdata(q_a_0),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_0),
	.prn(vcc));
defparam \MonDReg[0] .is_wysiwyg = "true";
defparam \MonDReg[0] .power_up = "low";

dffeas \MonDReg[24] (
	.clk(clk_clk),
	.d(jdo_27),
	.asdata(q_a_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_24),
	.prn(vcc));
defparam \MonDReg[24] .is_wysiwyg = "true";
defparam \MonDReg[24] .power_up = "low";

dffeas \MonDReg[4] (
	.clk(clk_clk),
	.d(jdo_7),
	.asdata(q_a_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_4),
	.prn(vcc));
defparam \MonDReg[4] .is_wysiwyg = "true";
defparam \MonDReg[4] .power_up = "low";

dffeas \MonDReg[20] (
	.clk(clk_clk),
	.d(jdo_23),
	.asdata(q_a_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_20),
	.prn(vcc));
defparam \MonDReg[20] .is_wysiwyg = "true";
defparam \MonDReg[20] .power_up = "low";

dffeas \MonDReg[19] (
	.clk(clk_clk),
	.d(jdo_22),
	.asdata(q_a_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_19),
	.prn(vcc));
defparam \MonDReg[19] .is_wysiwyg = "true";
defparam \MonDReg[19] .power_up = "low";

dffeas \MonDReg[16] (
	.clk(clk_clk),
	.d(jdo_19),
	.asdata(q_a_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_16),
	.prn(vcc));
defparam \MonDReg[16] .is_wysiwyg = "true";
defparam \MonDReg[16] .power_up = "low";

dffeas \MonDReg[25] (
	.clk(clk_clk),
	.d(jdo_28),
	.asdata(q_a_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_25),
	.prn(vcc));
defparam \MonDReg[25] .is_wysiwyg = "true";
defparam \MonDReg[25] .power_up = "low";

dffeas \MonDReg[26] (
	.clk(clk_clk),
	.d(jdo_29),
	.asdata(q_a_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_26),
	.prn(vcc));
defparam \MonDReg[26] .is_wysiwyg = "true";
defparam \MonDReg[26] .power_up = "low";

dffeas \MonDReg[27] (
	.clk(clk_clk),
	.d(jdo_30),
	.asdata(q_a_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_27),
	.prn(vcc));
defparam \MonDReg[27] .is_wysiwyg = "true";
defparam \MonDReg[27] .power_up = "low";

dffeas \MonDReg[28] (
	.clk(clk_clk),
	.d(jdo_31),
	.asdata(q_a_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_28),
	.prn(vcc));
defparam \MonDReg[28] .is_wysiwyg = "true";
defparam \MonDReg[28] .power_up = "low";

dffeas \MonDReg[30] (
	.clk(clk_clk),
	.d(jdo_33),
	.asdata(q_a_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_30),
	.prn(vcc));
defparam \MonDReg[30] .is_wysiwyg = "true";
defparam \MonDReg[30] .power_up = "low";

dffeas \MonDReg[31] (
	.clk(clk_clk),
	.d(jdo_34),
	.asdata(q_a_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_31),
	.prn(vcc));
defparam \MonDReg[31] .is_wysiwyg = "true";
defparam \MonDReg[31] .power_up = "low";

dffeas \MonDReg[21] (
	.clk(clk_clk),
	.d(jdo_24),
	.asdata(q_a_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_21),
	.prn(vcc));
defparam \MonDReg[21] .is_wysiwyg = "true";
defparam \MonDReg[21] .power_up = "low";

dffeas \MonDReg[17] (
	.clk(clk_clk),
	.d(jdo_20),
	.asdata(q_a_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_17),
	.prn(vcc));
defparam \MonDReg[17] .is_wysiwyg = "true";
defparam \MonDReg[17] .power_up = "low";

dffeas \MonDReg[6] (
	.clk(clk_clk),
	.d(jdo_9),
	.asdata(q_a_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_6),
	.prn(vcc));
defparam \MonDReg[6] .is_wysiwyg = "true";
defparam \MonDReg[6] .power_up = "low";

dffeas \MonDReg[22] (
	.clk(clk_clk),
	.d(jdo_25),
	.asdata(q_a_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_22),
	.prn(vcc));
defparam \MonDReg[22] .is_wysiwyg = "true";
defparam \MonDReg[22] .power_up = "low";

dffeas \MonDReg[23] (
	.clk(clk_clk),
	.d(jdo_26),
	.asdata(q_a_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_23),
	.prn(vcc));
defparam \MonDReg[23] .is_wysiwyg = "true";
defparam \MonDReg[23] .power_up = "low";

dffeas \MonDReg[7] (
	.clk(clk_clk),
	.d(jdo_10),
	.asdata(q_a_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_7),
	.prn(vcc));
defparam \MonDReg[7] .is_wysiwyg = "true";
defparam \MonDReg[7] .power_up = "low";

dffeas \MonDReg[15] (
	.clk(clk_clk),
	.d(jdo_18),
	.asdata(q_a_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_15),
	.prn(vcc));
defparam \MonDReg[15] .is_wysiwyg = "true";
defparam \MonDReg[15] .power_up = "low";

dffeas \MonDReg[13] (
	.clk(clk_clk),
	.d(jdo_16),
	.asdata(q_a_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_13),
	.prn(vcc));
defparam \MonDReg[13] .is_wysiwyg = "true";
defparam \MonDReg[13] .power_up = "low";

dffeas \MonDReg[14] (
	.clk(clk_clk),
	.d(jdo_17),
	.asdata(q_a_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\MonDReg[23]~0_combout ),
	.sload(!take_action_ocimem_b),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_14),
	.prn(vcc));
defparam \MonDReg[14] .is_wysiwyg = "true";
defparam \MonDReg[14] .power_up = "low";

dffeas waitrequest(
	.clk(clk_clk),
	.d(\waitrequest~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(waitrequest1),
	.prn(vcc));
defparam waitrequest.is_wysiwyg = "true";
defparam waitrequest.power_up = "low";

dffeas \MonDReg[1] (
	.clk(clk_clk),
	.d(\MonDReg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_1),
	.prn(vcc));
defparam \MonDReg[1] .is_wysiwyg = "true";
defparam \MonDReg[1] .power_up = "low";

dffeas \MonDReg[2] (
	.clk(clk_clk),
	.d(\MonDReg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_2),
	.prn(vcc));
defparam \MonDReg[2] .is_wysiwyg = "true";
defparam \MonDReg[2] .power_up = "low";

dffeas \MonDReg[3] (
	.clk(clk_clk),
	.d(\MonDReg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_3),
	.prn(vcc));
defparam \MonDReg[3] .is_wysiwyg = "true";
defparam \MonDReg[3] .power_up = "low";

dffeas \MonDReg[5] (
	.clk(clk_clk),
	.d(\MonDReg~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_5),
	.prn(vcc));
defparam \MonDReg[5] .is_wysiwyg = "true";
defparam \MonDReg[5] .power_up = "low";

dffeas \MonDReg[29] (
	.clk(clk_clk),
	.d(\MonDReg~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_29),
	.prn(vcc));
defparam \MonDReg[29] .is_wysiwyg = "true";
defparam \MonDReg[29] .power_up = "low";

dffeas \MonDReg[18] (
	.clk(clk_clk),
	.d(\MonDReg~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_18),
	.prn(vcc));
defparam \MonDReg[18] .is_wysiwyg = "true";
defparam \MonDReg[18] .power_up = "low";

dffeas \MonDReg[10] (
	.clk(clk_clk),
	.d(\MonDReg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_10),
	.prn(vcc));
defparam \MonDReg[10] .is_wysiwyg = "true";
defparam \MonDReg[10] .power_up = "low";

dffeas \MonDReg[12] (
	.clk(clk_clk),
	.d(\MonDReg[12]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[12]~8_combout ),
	.q(MonDReg_12),
	.prn(vcc));
defparam \MonDReg[12] .is_wysiwyg = "true";
defparam \MonDReg[12] .power_up = "low";

dffeas \MonDReg[11] (
	.clk(clk_clk),
	.d(\MonDReg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_11),
	.prn(vcc));
defparam \MonDReg[11] .is_wysiwyg = "true";
defparam \MonDReg[11] .power_up = "low";

dffeas \MonDReg[9] (
	.clk(clk_clk),
	.d(\MonDReg~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[0]~1_combout ),
	.q(MonDReg_9),
	.prn(vcc));
defparam \MonDReg[9] .is_wysiwyg = "true";
defparam \MonDReg[9] .power_up = "low";

dffeas \MonDReg[8] (
	.clk(clk_clk),
	.d(\MonDReg[8]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\MonDReg[12]~8_combout ),
	.q(MonDReg_8),
	.prn(vcc));
defparam \MonDReg[8] .is_wysiwyg = "true";
defparam \MonDReg[8] .power_up = "low";

cyclonev_lcell_comb \Add0~1_wirecell (
	.dataa(!\Add0~1_sumout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_wirecell_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1_wirecell .extended_lut = "off";
defparam \Add0~1_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \Add0~1_wirecell .shared_arith = "off";

dffeas \MonAReg[10] (
	.clk(clk_clk),
	.d(\Add0~1_wirecell_combout ),
	.asdata(jdo_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[10]~q ),
	.prn(vcc));
defparam \MonAReg[10] .is_wysiwyg = "true";
defparam \MonAReg[10] .power_up = "low";

cyclonev_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[2]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \MonAReg[2] (
	.clk(clk_clk),
	.d(\Add0~9_sumout ),
	.asdata(jdo_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[2]~q ),
	.prn(vcc));
defparam \MonAReg[2] .is_wysiwyg = "true";
defparam \MonAReg[2] .power_up = "low";

cyclonev_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \MonAReg[3] (
	.clk(clk_clk),
	.d(\Add0~5_sumout ),
	.asdata(jdo_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[3]~q ),
	.prn(vcc));
defparam \MonAReg[3] .is_wysiwyg = "true";
defparam \MonAReg[3] .power_up = "low";

cyclonev_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \MonAReg[4] (
	.clk(clk_clk),
	.d(\Add0~13_sumout ),
	.asdata(jdo_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[4]~q ),
	.prn(vcc));
defparam \MonAReg[4] .is_wysiwyg = "true";
defparam \MonAReg[4] .power_up = "low";

cyclonev_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[5]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \MonAReg[5] (
	.clk(clk_clk),
	.d(\Add0~17_sumout ),
	.asdata(jdo_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[5]~q ),
	.prn(vcc));
defparam \MonAReg[5] .is_wysiwyg = "true";
defparam \MonAReg[5] .power_up = "low";

cyclonev_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[6]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \MonAReg[6] (
	.clk(clk_clk),
	.d(\Add0~21_sumout ),
	.asdata(jdo_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[6]~q ),
	.prn(vcc));
defparam \MonAReg[6] .is_wysiwyg = "true";
defparam \MonAReg[6] .power_up = "low";

cyclonev_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[7]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \MonAReg[7] (
	.clk(clk_clk),
	.d(\Add0~25_sumout ),
	.asdata(jdo_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[7]~q ),
	.prn(vcc));
defparam \MonAReg[7] .is_wysiwyg = "true";
defparam \MonAReg[7] .power_up = "low";

cyclonev_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[8]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \MonAReg[8] (
	.clk(clk_clk),
	.d(\Add0~29_sumout ),
	.asdata(jdo_32),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[8]~q ),
	.prn(vcc));
defparam \MonAReg[8] .is_wysiwyg = "true";
defparam \MonAReg[8] .power_up = "low";

cyclonev_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \MonAReg[9] (
	.clk(clk_clk),
	.d(\Add0~33_sumout ),
	.asdata(jdo_33),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(take_action_ocimem_a2),
	.ena(take_action_ocimem_a),
	.q(\MonAReg[9]~q ),
	.prn(vcc));
defparam \MonAReg[9] .is_wysiwyg = "true";
defparam \MonAReg[9] .power_up = "low";

cyclonev_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\MonAReg[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_rd~0 (
	.dataa(!take_action_ocimem_a1),
	.datab(!jdo_34),
	.datac(!jdo_17),
	.datad(!\Add0~1_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_rd~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_rd~0 .extended_lut = "off";
defparam \jtag_ram_rd~0 .lut_mask = 64'hD1FFD1FFD1FFD1FF;
defparam \jtag_ram_rd~0 .shared_arith = "off";

dffeas jtag_ram_rd(
	.clk(clk_clk),
	.d(\jtag_ram_rd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_action_ocimem_b),
	.q(\jtag_ram_rd~q ),
	.prn(vcc));
defparam jtag_ram_rd.is_wysiwyg = "true";
defparam jtag_ram_rd.power_up = "low";

dffeas jtag_ram_rd_d1(
	.clk(clk_clk),
	.d(\jtag_ram_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_rd_d1~q ),
	.prn(vcc));
defparam jtag_ram_rd_d1.is_wysiwyg = "true";
defparam jtag_ram_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[23]~0 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!take_action_ocimem_b),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[23]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[23]~0 .extended_lut = "off";
defparam \MonDReg[23]~0 .lut_mask = 64'hEEEEEEEEEEEEEEEE;
defparam \MonDReg[23]~0 .shared_arith = "off";

dffeas jtag_rd(
	.clk(clk_clk),
	.d(take_action_ocimem_a1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(!take_action_ocimem_b),
	.q(\jtag_rd~q ),
	.prn(vcc));
defparam jtag_rd.is_wysiwyg = "true";
defparam jtag_rd.power_up = "low";

dffeas jtag_rd_d1(
	.clk(clk_clk),
	.d(\jtag_rd~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_rd_d1~q ),
	.prn(vcc));
defparam jtag_rd_d1.is_wysiwyg = "true";
defparam jtag_rd_d1.power_up = "low";

cyclonev_lcell_comb \MonDReg[0]~1 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_35),
	.datac(!\jtag_rd_d1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[0]~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[0]~1 .extended_lut = "off";
defparam \MonDReg[0]~1 .lut_mask = 64'h2727272727272727;
defparam \MonDReg[0]~1 .shared_arith = "off";

cyclonev_lcell_comb \jtag_ram_access~0 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_35),
	.datac(!jdo_34),
	.datad(!jdo_17),
	.datae(!\Add0~1_sumout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\jtag_ram_access~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \jtag_ram_access~0 .extended_lut = "off";
defparam \jtag_ram_access~0 .lut_mask = 64'hFF7DFFFFFF7DFFFF;
defparam \jtag_ram_access~0 .shared_arith = "off";

dffeas jtag_ram_access(
	.clk(clk_clk),
	.d(\jtag_ram_access~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\jtag_ram_access~q ),
	.prn(vcc));
defparam jtag_ram_access.is_wysiwyg = "true";
defparam jtag_ram_access.power_up = "low";

cyclonev_lcell_comb \waitrequest~0 (
	.dataa(!address_8),
	.datab(!\jtag_ram_access~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~0 .extended_lut = "off";
defparam \waitrequest~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \waitrequest~0 .shared_arith = "off";

cyclonev_lcell_comb \avalon_ociram_readdata_ready~0 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\avalon_ociram_readdata_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \avalon_ociram_readdata_ready~0 .extended_lut = "off";
defparam \avalon_ociram_readdata_ready~0 .lut_mask = 64'hD1FFFFFFD1FFFFFF;
defparam \avalon_ociram_readdata_ready~0 .shared_arith = "off";

dffeas avalon_ociram_readdata_ready(
	.clk(clk_clk),
	.d(\avalon_ociram_readdata_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\avalon_ociram_readdata_ready~q ),
	.prn(vcc));
defparam avalon_ociram_readdata_ready.is_wysiwyg = "true";
defparam avalon_ociram_readdata_ready.power_up = "low";

cyclonev_lcell_comb \waitrequest~1 (
	.dataa(!waitrequest1),
	.datab(!write),
	.datac(!\waitrequest~0_combout ),
	.datad(!read),
	.datae(!\avalon_ociram_readdata_ready~q ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\waitrequest~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \waitrequest~1 .extended_lut = "off";
defparam \waitrequest~1 .lut_mask = 64'hFFFFBF8FFFFFBF8F;
defparam \waitrequest~1 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~2 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[2]~q ),
	.datad(!\MonAReg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~2 .extended_lut = "off";
defparam \MonDReg~2 .lut_mask = 64'hFFEFFFEFFFEFFFEF;
defparam \MonDReg~2 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~3 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!take_action_ocimem_b),
	.datac(!jdo_4),
	.datad(!q_a_1),
	.datae(!\MonDReg~2_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~3 .extended_lut = "off";
defparam \MonDReg~3 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~3 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~4 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!\MonAReg[3]~q ),
	.datac(!\MonAReg[2]~q ),
	.datad(!\MonAReg[4]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~4 .extended_lut = "off";
defparam \MonDReg~4 .lut_mask = 64'hEFFEEFFEEFFEEFFE;
defparam \MonDReg~4 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~5 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!take_action_ocimem_b),
	.datac(!jdo_5),
	.datad(!q_a_2),
	.datae(!\MonDReg~4_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~5 .extended_lut = "off";
defparam \MonDReg~5 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~5 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~6 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!take_action_ocimem_b),
	.datac(!\MonDReg~4_combout ),
	.datad(!jdo_6),
	.datae(!q_a_3),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~6 .extended_lut = "off";
defparam \MonDReg~6 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~6 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~27 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!q_a_5),
	.datad(!jdo_8),
	.datae(!\jtag_ram_rd_d1~q ),
	.dataf(!take_action_ocimem_b),
	.datag(!\MonAReg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~27_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~27 .extended_lut = "on";
defparam \MonDReg~27 .lut_mask = 64'hFF7FFFF7FF7FFFF7;
defparam \MonDReg~27 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~23 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!q_a_29),
	.datad(!jdo_32),
	.datae(!\jtag_ram_rd_d1~q ),
	.dataf(!take_action_ocimem_b),
	.datag(!\MonAReg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~23_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~23 .extended_lut = "on";
defparam \MonDReg~23 .lut_mask = 64'hFFBFFFFBFFBFFFFB;
defparam \MonDReg~23 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~19 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!q_a_18),
	.datad(!jdo_21),
	.datae(!\jtag_ram_rd_d1~q ),
	.dataf(!take_action_ocimem_b),
	.datag(!\MonAReg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~19_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~19 .extended_lut = "on";
defparam \MonDReg~19 .lut_mask = 64'hFFF7FFF7FFF7FFF7;
defparam \MonDReg~19 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~7 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!take_action_ocimem_b),
	.datac(!\MonDReg~2_combout ),
	.datad(!q_a_10),
	.datae(!jdo_13),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~7 .extended_lut = "off";
defparam \MonDReg~7 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~7 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[12]~15 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!q_a_12),
	.datad(!jdo_15),
	.datae(!\jtag_ram_rd_d1~q ),
	.dataf(!take_action_ocimem_b),
	.datag(!\MonAReg[3]~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[12]~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[12]~15 .extended_lut = "on";
defparam \MonDReg[12]~15 .lut_mask = 64'hFF6FFFF6FF6FFFF6;
defparam \MonDReg[12]~15 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[12]~8 (
	.dataa(!take_action_ocimem_a),
	.datab(!jdo_35),
	.datac(!\jtag_rd_d1~q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[12]~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[12]~8 .extended_lut = "off";
defparam \MonDReg[12]~8 .lut_mask = 64'h2727272727272727;
defparam \MonDReg[12]~8 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~9 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!take_action_ocimem_b),
	.datac(!\MonDReg~4_combout ),
	.datad(!q_a_11),
	.datae(!jdo_14),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~9 .extended_lut = "off";
defparam \MonDReg~9 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~9 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg~10 (
	.dataa(!\jtag_ram_rd_d1~q ),
	.datab(!take_action_ocimem_b),
	.datac(!\MonDReg~4_combout ),
	.datad(!q_a_9),
	.datae(!jdo_12),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg~10 .extended_lut = "off";
defparam \MonDReg~10 .lut_mask = 64'h47FFFFFF47FFFFFF;
defparam \MonDReg~10 .shared_arith = "off";

cyclonev_lcell_comb \MonDReg[8]~11 (
	.dataa(!\MonAReg[4]~q ),
	.datab(!\MonAReg[2]~q ),
	.datac(!jdo_11),
	.datad(!\MonAReg[3]~q ),
	.datae(!take_action_ocimem_b),
	.dataf(!q_a_8),
	.datag(!\jtag_ram_rd_d1~q ),
	.cin(gnd),
	.sharein(gnd),
	.combout(\MonDReg[8]~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \MonDReg[8]~11 .extended_lut = "on";
defparam \MonDReg[8]~11 .lut_mask = 64'h6996F9F66996F9F6;
defparam \MonDReg[8]~11 .shared_arith = "off";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_ociram_sp_ram_module (
	q_a_0,
	q_a_1,
	q_a_2,
	q_a_3,
	q_a_24,
	q_a_4,
	q_a_20,
	q_a_19,
	q_a_16,
	q_a_25,
	q_a_5,
	q_a_26,
	q_a_27,
	q_a_28,
	q_a_29,
	q_a_30,
	q_a_31,
	q_a_21,
	q_a_18,
	q_a_17,
	q_a_10,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_13,
	q_a_12,
	q_a_11,
	q_a_9,
	q_a_8,
	q_a_6,
	q_a_14,
	q_a_22,
	ociram_wr_en,
	ociram_reset_req,
	ociram_wr_data_0,
	ociram_addr_0,
	ociram_addr_1,
	ociram_addr_2,
	ociram_addr_3,
	ociram_addr_4,
	ociram_addr_5,
	ociram_addr_6,
	ociram_addr_7,
	ociram_byteenable_0,
	ociram_wr_data_1,
	ociram_wr_data_2,
	ociram_wr_data_3,
	ociram_wr_data_24,
	ociram_byteenable_3,
	ociram_wr_data_4,
	ociram_wr_data_20,
	ociram_byteenable_2,
	ociram_wr_data_19,
	ociram_wr_data_16,
	ociram_wr_data_25,
	ociram_wr_data_5,
	ociram_wr_data_26,
	ociram_wr_data_27,
	ociram_wr_data_28,
	ociram_wr_data_29,
	ociram_wr_data_30,
	ociram_wr_data_31,
	ociram_wr_data_21,
	ociram_wr_data_18,
	ociram_wr_data_17,
	ociram_wr_data_10,
	ociram_byteenable_1,
	ociram_wr_data_7,
	ociram_wr_data_23,
	ociram_wr_data_15,
	ociram_wr_data_13,
	ociram_wr_data_12,
	ociram_wr_data_11,
	ociram_wr_data_9,
	ociram_wr_data_8,
	ociram_wr_data_6,
	ociram_wr_data_14,
	ociram_wr_data_22,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_a_1;
output 	q_a_2;
output 	q_a_3;
output 	q_a_24;
output 	q_a_4;
output 	q_a_20;
output 	q_a_19;
output 	q_a_16;
output 	q_a_25;
output 	q_a_5;
output 	q_a_26;
output 	q_a_27;
output 	q_a_28;
output 	q_a_29;
output 	q_a_30;
output 	q_a_31;
output 	q_a_21;
output 	q_a_18;
output 	q_a_17;
output 	q_a_10;
output 	q_a_7;
output 	q_a_23;
output 	q_a_15;
output 	q_a_13;
output 	q_a_12;
output 	q_a_11;
output 	q_a_9;
output 	q_a_8;
output 	q_a_6;
output 	q_a_14;
output 	q_a_22;
input 	ociram_wr_en;
input 	ociram_reset_req;
input 	ociram_wr_data_0;
input 	ociram_addr_0;
input 	ociram_addr_1;
input 	ociram_addr_2;
input 	ociram_addr_3;
input 	ociram_addr_4;
input 	ociram_addr_5;
input 	ociram_addr_6;
input 	ociram_addr_7;
input 	ociram_byteenable_0;
input 	ociram_wr_data_1;
input 	ociram_wr_data_2;
input 	ociram_wr_data_3;
input 	ociram_wr_data_24;
input 	ociram_byteenable_3;
input 	ociram_wr_data_4;
input 	ociram_wr_data_20;
input 	ociram_byteenable_2;
input 	ociram_wr_data_19;
input 	ociram_wr_data_16;
input 	ociram_wr_data_25;
input 	ociram_wr_data_5;
input 	ociram_wr_data_26;
input 	ociram_wr_data_27;
input 	ociram_wr_data_28;
input 	ociram_wr_data_29;
input 	ociram_wr_data_30;
input 	ociram_wr_data_31;
input 	ociram_wr_data_21;
input 	ociram_wr_data_18;
input 	ociram_wr_data_17;
input 	ociram_wr_data_10;
input 	ociram_byteenable_1;
input 	ociram_wr_data_7;
input 	ociram_wr_data_23;
input 	ociram_wr_data_15;
input 	ociram_wr_data_13;
input 	ociram_wr_data_12;
input 	ociram_wr_data_11;
input 	ociram_wr_data_9;
input 	ociram_wr_data_8;
input 	ociram_wr_data_6;
input 	ociram_wr_data_14;
input 	ociram_wr_data_22;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_7 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.wren_a(ociram_wr_en),
	.clocken0(ociram_reset_req),
	.data_a({ociram_wr_data_31,ociram_wr_data_30,ociram_wr_data_29,ociram_wr_data_28,ociram_wr_data_27,ociram_wr_data_26,ociram_wr_data_25,ociram_wr_data_24,ociram_wr_data_23,ociram_wr_data_22,ociram_wr_data_21,ociram_wr_data_20,ociram_wr_data_19,ociram_wr_data_18,ociram_wr_data_17,
ociram_wr_data_16,ociram_wr_data_15,ociram_wr_data_14,ociram_wr_data_13,ociram_wr_data_12,ociram_wr_data_11,ociram_wr_data_10,ociram_wr_data_9,ociram_wr_data_8,ociram_wr_data_7,ociram_wr_data_6,ociram_wr_data_5,ociram_wr_data_4,ociram_wr_data_3,ociram_wr_data_2,
ociram_wr_data_1,ociram_wr_data_0}),
	.address_a({gnd,gnd,ociram_addr_7,ociram_addr_6,ociram_addr_5,ociram_addr_4,ociram_addr_3,ociram_addr_2,ociram_addr_1,ociram_addr_0}),
	.byteena_a({ociram_byteenable_3,ociram_byteenable_2,ociram_byteenable_1,ociram_byteenable_0}),
	.clock0(clk_clk));

endmodule

module embedded_system_altsyncram_7 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[9:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_j7g1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.wren_a(wren_a),
	.clocken0(clocken0),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module embedded_system_altsyncram_j7g1 (
	q_a,
	wren_a,
	clocken0,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	wren_a;
input 	clocken0;
input 	[31:0] data_a;
input 	[7:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 8;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 255;
defparam ram_block1a0.port_a_logical_ram_depth = 256;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "2080506BCF0D06D1F082E980277062912CB244CFD084FC8EC49C6B4F28A56006";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 8;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 255;
defparam ram_block1a1.port_a_logical_ram_depth = 256;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "66F9986418FBBDC2D79799D62A2EBCDE87554821870A4291446385CAE645D15F";

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 8;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 255;
defparam ram_block1a2.port_a_logical_ram_depth = 256;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "633A992C2A4C071E706E6722D5D1FDC707F573CF0D406D54B651FC97C911E5D3";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 8;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 255;
defparam ram_block1a3.port_a_logical_ram_depth = 256;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "4F950EEE46E51336E633C4C82AD564200DDC93F4E4FCFE0F10D3E8843064AB49";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 8;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 255;
defparam ram_block1a24.port_a_logical_ram_depth = 256;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = "1611CFF2626AB6D5471DD74C4854A7C640358F5D02EF6605C204E43D41486417";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 8;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 255;
defparam ram_block1a4.port_a_logical_ram_depth = 256;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "0C89DA0AC7212C6B79E89849B2238B9BB6E73FE43D9BC8C166A1F9C0F6BA1EAA";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 8;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 255;
defparam ram_block1a20.port_a_logical_ram_depth = 256;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "4C0DBABA3E5B0DC65CF4DC015DC4B93CAC73E3F541C878BD0279B1FC525FA32A";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 8;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 255;
defparam ram_block1a19.port_a_logical_ram_depth = 256;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "8BB0528D733F0CE7360DDF4DBED01AA957F9DF48CA69E672F9EEDAFEAC738A5C";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 8;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 255;
defparam ram_block1a16.port_a_logical_ram_depth = 256;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "D3BF8815D6EA52ACA5D90182D0FEE54279153DC162279DA35E59C350C65ACE27";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 8;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 255;
defparam ram_block1a25.port_a_logical_ram_depth = 256;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = "6047012728D997AD87894BF09AAB5618DC7D301FAFF1AB6CCC1AFF1791A2DF6D";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 8;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 255;
defparam ram_block1a5.port_a_logical_ram_depth = 256;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "B9B1E2FF67F9B8C056385C7763CD70C3C6A16547526E3BE75D897A6DE98AB7B6";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 8;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 255;
defparam ram_block1a26.port_a_logical_ram_depth = 256;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = "737C19A08111F0CD2B4C4C58C3FB8AF5BED936D1221A104CAA70AAD527639343";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 8;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 255;
defparam ram_block1a27.port_a_logical_ram_depth = 256;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = "0B3AE958620CF874FB552A1D483607D3E50925BCD213C99CC386063369FA8A9C";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 8;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 255;
defparam ram_block1a28.port_a_logical_ram_depth = 256;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = "D2FACB3874CB7F69A2230993CF91AB682BECD42F86F5803561257952176173A7";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 8;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 255;
defparam ram_block1a29.port_a_logical_ram_depth = 256;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = "9F4ED31DC21880DB480F616A1CF268494538501BEFD54167C5679AB6979341F9";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 8;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 255;
defparam ram_block1a30.port_a_logical_ram_depth = 256;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = "F5641D6C8836BF000D1DCE468A1830B27E519D02FAF7E48644C58296B6B82905";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 8;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 255;
defparam ram_block1a31.port_a_logical_ram_depth = 256;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = "6508DD5113A38E018C39BEA8FC3C6D2B053FC6729A29ACA3A834D004F11037B3";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 8;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 255;
defparam ram_block1a21.port_a_logical_ram_depth = 256;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "B0CD28E8539066BFB50B0604E542D1D67047F6548C867D78F987A48D04D1CA5C";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 8;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 255;
defparam ram_block1a18.port_a_logical_ram_depth = 256;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "9EDD4BC3F1041988DEF2B79C2B0A6D738AD7EB2EFDC138C31CA5C1478DB6AE9D";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 8;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 255;
defparam ram_block1a17.port_a_logical_ram_depth = 256;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "90F92BF4047F2973C1F7B73EE93A06E9824DC9DAEC9FDFADDB2ACDCFC8DEFA54";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 8;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 255;
defparam ram_block1a10.port_a_logical_ram_depth = 256;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "ABBA72442BE0093687C0D5782816FE7CE5847E0EC072EE77BF6263BECDFF886C";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 8;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 255;
defparam ram_block1a7.port_a_logical_ram_depth = 256;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "9E4C1F6675D4244D809042A238CD1915199CC77B204E9890128E2108FD03AF3C";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 8;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 255;
defparam ram_block1a23.port_a_logical_ram_depth = 256;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "04BE6ABADBE8C2C2F2FF32884A75FB4E414BCC5ED0D90F02E051607E45864981";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 8;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 255;
defparam ram_block1a15.port_a_logical_ram_depth = 256;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "56BE0FCB022E30A1E454C43F0A08EDEA0EE78B116A19AFE6DB876AD24EC24281";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 8;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 255;
defparam ram_block1a13.port_a_logical_ram_depth = 256;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "8105F14E5EEC9F1AD891C645AC0EC442B741340091FA518E10D334A5CC003D79";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 8;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 255;
defparam ram_block1a12.port_a_logical_ram_depth = 256;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "13F7E86ED8B5C2E0CAFE8146F9752B2065A8CED2B02561410CA1B76131DB11AC";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 8;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 255;
defparam ram_block1a11.port_a_logical_ram_depth = 256;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "A8A81B1AAAD3D7D688E515FCA96491A7760B8047458582F91DAF2659A83C0CB0";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 8;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 255;
defparam ram_block1a9.port_a_logical_ram_depth = 256;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "62A2C8A25E376C028612C41166A7972AFBFFC4A72AA1DEC34D8048511E87B0B1";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 8;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 255;
defparam ram_block1a8.port_a_logical_ram_depth = 256;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "5E8E2CCA3F98B355B4D77C1E3C88B38DC941C69776E33B1C652A6C84E8833864";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 8;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 255;
defparam ram_block1a6.port_a_logical_ram_depth = 256;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "F0BA9F8E9501E35ED88C8AC651B0172375610EAA646E019096C91D55B564B1D3";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 8;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 255;
defparam ram_block1a14.port_a_logical_ram_depth = 256;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "C6A4915740F2841D3E15CCDE46521E7FCEBD107E14CF06B37D5ED68D563B69BD";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "embedded_system_nios2_qsys_0_ociram_default_contents.mif";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_nios2_oci:the_embedded_system_nios2_qsys_0_nios2_oci|embedded_system_nios2_qsys_0_nios2_ocimem:the_embedded_system_nios2_qsys_0_nios2_ocimem|embedded_system_nios2_qsys_0_ociram_sp_ram_module:embedded_system_nios2_qsys_0_ociram_sp_ram|altsyncram:the_altsyncram|altsyncram_j7g1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 8;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 255;
defparam ram_block1a22.port_a_logical_ram_depth = 256;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "5FF25143060CBCF9A3D3B17971E078A0354875B91E2AA9D03DE4032006CE8686";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_register_bank_a_module (
	q_b_2,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_27,
	q_b_29,
	q_b_30,
	q_b_31,
	q_b_17,
	q_b_16,
	q_b_28,
	q_b_18,
	q_b_26,
	q_b_19,
	q_b_21,
	q_b_15,
	q_b_25,
	q_b_20,
	q_b_22,
	q_b_14,
	q_b_24,
	q_b_23,
	q_b_1,
	q_b_0,
	A_wr_data_unfiltered_2,
	A_wr_data_unfiltered_13,
	A_wr_data_unfiltered_12,
	A_wr_data_unfiltered_11,
	A_wr_data_unfiltered_10,
	A_wr_data_unfiltered_9,
	A_wr_data_unfiltered_8,
	A_wr_data_unfiltered_7,
	A_wr_data_unfiltered_6,
	A_wr_data_unfiltered_5,
	A_wr_data_unfiltered_4,
	A_wr_data_unfiltered_3,
	A_wr_data_unfiltered_1,
	A_wr_data_unfiltered_0,
	A_wr_data_unfiltered_21,
	A_wr_data_unfiltered_20,
	A_wr_data_unfiltered_25,
	A_wr_data_unfiltered_17,
	A_wr_data_unfiltered_24,
	A_wr_data_unfiltered_16,
	A_wr_data_unfiltered_27,
	A_wr_data_unfiltered_19,
	A_wr_data_unfiltered_26,
	A_wr_data_unfiltered_18,
	A_wr_data_unfiltered_23,
	A_wr_data_unfiltered_22,
	A_wr_data_unfiltered_29,
	A_wr_data_unfiltered_30,
	A_wr_data_unfiltered_31,
	A_wr_data_unfiltered_28,
	A_wr_data_unfiltered_15,
	A_wr_data_unfiltered_14,
	A_dst_regnum_from_M_4,
	A_wr_dst_reg_from_M,
	A_dst_regnum_from_M_0,
	A_dst_regnum_from_M_1,
	A_dst_regnum_from_M_2,
	A_dst_regnum_from_M_3,
	rf_a_rd_port_addr_0,
	rf_a_rd_port_addr_1,
	rf_a_rd_port_addr_2,
	rf_a_rd_port_addr_3,
	rf_a_rd_port_addr_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_2;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_27;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
output 	q_b_17;
output 	q_b_16;
output 	q_b_28;
output 	q_b_18;
output 	q_b_26;
output 	q_b_19;
output 	q_b_21;
output 	q_b_15;
output 	q_b_25;
output 	q_b_20;
output 	q_b_22;
output 	q_b_14;
output 	q_b_24;
output 	q_b_23;
output 	q_b_1;
output 	q_b_0;
input 	A_wr_data_unfiltered_2;
input 	A_wr_data_unfiltered_13;
input 	A_wr_data_unfiltered_12;
input 	A_wr_data_unfiltered_11;
input 	A_wr_data_unfiltered_10;
input 	A_wr_data_unfiltered_9;
input 	A_wr_data_unfiltered_8;
input 	A_wr_data_unfiltered_7;
input 	A_wr_data_unfiltered_6;
input 	A_wr_data_unfiltered_5;
input 	A_wr_data_unfiltered_4;
input 	A_wr_data_unfiltered_3;
input 	A_wr_data_unfiltered_1;
input 	A_wr_data_unfiltered_0;
input 	A_wr_data_unfiltered_21;
input 	A_wr_data_unfiltered_20;
input 	A_wr_data_unfiltered_25;
input 	A_wr_data_unfiltered_17;
input 	A_wr_data_unfiltered_24;
input 	A_wr_data_unfiltered_16;
input 	A_wr_data_unfiltered_27;
input 	A_wr_data_unfiltered_19;
input 	A_wr_data_unfiltered_26;
input 	A_wr_data_unfiltered_18;
input 	A_wr_data_unfiltered_23;
input 	A_wr_data_unfiltered_22;
input 	A_wr_data_unfiltered_29;
input 	A_wr_data_unfiltered_30;
input 	A_wr_data_unfiltered_31;
input 	A_wr_data_unfiltered_28;
input 	A_wr_data_unfiltered_15;
input 	A_wr_data_unfiltered_14;
input 	A_dst_regnum_from_M_4;
input 	A_wr_dst_reg_from_M;
input 	A_dst_regnum_from_M_0;
input 	A_dst_regnum_from_M_1;
input 	A_dst_regnum_from_M_2;
input 	A_dst_regnum_from_M_3;
input 	rf_a_rd_port_addr_0;
input 	rf_a_rd_port_addr_1;
input 	rf_a_rd_port_addr_2;
input 	rf_a_rd_port_addr_3;
input 	rf_a_rd_port_addr_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_8 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({A_wr_data_unfiltered_31,A_wr_data_unfiltered_30,A_wr_data_unfiltered_29,A_wr_data_unfiltered_28,A_wr_data_unfiltered_27,A_wr_data_unfiltered_26,A_wr_data_unfiltered_25,A_wr_data_unfiltered_24,A_wr_data_unfiltered_23,A_wr_data_unfiltered_22,A_wr_data_unfiltered_21,
A_wr_data_unfiltered_20,A_wr_data_unfiltered_19,A_wr_data_unfiltered_18,A_wr_data_unfiltered_17,A_wr_data_unfiltered_16,A_wr_data_unfiltered_15,A_wr_data_unfiltered_14,A_wr_data_unfiltered_13,A_wr_data_unfiltered_12,A_wr_data_unfiltered_11,A_wr_data_unfiltered_10,
A_wr_data_unfiltered_9,A_wr_data_unfiltered_8,A_wr_data_unfiltered_7,A_wr_data_unfiltered_6,A_wr_data_unfiltered_5,A_wr_data_unfiltered_4,A_wr_data_unfiltered_3,A_wr_data_unfiltered_2,A_wr_data_unfiltered_1,A_wr_data_unfiltered_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,A_dst_regnum_from_M_4,A_dst_regnum_from_M_3,A_dst_regnum_from_M_2,A_dst_regnum_from_M_1,A_dst_regnum_from_M_0}),
	.wren_a(A_wr_dst_reg_from_M),
	.address_b({gnd,gnd,gnd,gnd,gnd,rf_a_rd_port_addr_4,rf_a_rd_port_addr_3,rf_a_rd_port_addr_2,rf_a_rd_port_addr_1,rf_a_rd_port_addr_0}),
	.clock0(clk_clk));

endmodule

module embedded_system_altsyncram_8 (
	q_b,
	data_a,
	address_a,
	wren_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	[9:0] address_a;
input 	wren_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_9tn1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.wren_a(wren_a),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module embedded_system_altsyncram_9tn1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a13.init_file_layout = "port_b";
defparam ram_block1a13.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a12.init_file_layout = "port_b";
defparam ram_block1a12.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a11.init_file_layout = "port_b";
defparam ram_block1a11.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a10.init_file_layout = "port_b";
defparam ram_block1a10.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a9.init_file_layout = "port_b";
defparam ram_block1a9.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a8.init_file_layout = "port_b";
defparam ram_block1a8.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a7.init_file_layout = "port_b";
defparam ram_block1a7.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a6.init_file_layout = "port_b";
defparam ram_block1a6.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a5.init_file_layout = "port_b";
defparam ram_block1a5.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a27.init_file_layout = "port_b";
defparam ram_block1a27.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a29.init_file_layout = "port_b";
defparam ram_block1a29.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a30.init_file_layout = "port_b";
defparam ram_block1a30.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a31.init_file_layout = "port_b";
defparam ram_block1a31.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a17.init_file_layout = "port_b";
defparam ram_block1a17.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a16.init_file_layout = "port_b";
defparam ram_block1a16.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a28.init_file_layout = "port_b";
defparam ram_block1a28.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a18.init_file_layout = "port_b";
defparam ram_block1a18.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a26.init_file_layout = "port_b";
defparam ram_block1a26.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a19.init_file_layout = "port_b";
defparam ram_block1a19.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a21.init_file_layout = "port_b";
defparam ram_block1a21.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a15.init_file_layout = "port_b";
defparam ram_block1a15.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a25.init_file_layout = "port_b";
defparam ram_block1a25.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a20.init_file_layout = "port_b";
defparam ram_block1a20.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a22.init_file_layout = "port_b";
defparam ram_block1a22.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a14.init_file_layout = "port_b";
defparam ram_block1a14.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a24.init_file_layout = "port_b";
defparam ram_block1a24.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a23.init_file_layout = "port_b";
defparam ram_block1a23.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "embedded_system_nios2_qsys_0_rf_ram_a.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_a_module:embedded_system_nios2_qsys_0_register_bank_a|altsyncram:the_altsyncram|altsyncram_9tn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "FFFFFFFF";

endmodule

module embedded_system_embedded_system_nios2_qsys_0_register_bank_b_module (
	q_b_2,
	q_b_13,
	q_b_12,
	q_b_11,
	q_b_10,
	q_b_9,
	q_b_8,
	q_b_7,
	q_b_6,
	q_b_5,
	q_b_4,
	q_b_3,
	q_b_1,
	q_b_0,
	q_b_21,
	q_b_20,
	q_b_25,
	q_b_17,
	q_b_24,
	q_b_16,
	q_b_27,
	q_b_19,
	q_b_26,
	q_b_18,
	q_b_23,
	q_b_15,
	q_b_22,
	q_b_14,
	q_b_29,
	q_b_30,
	q_b_31,
	q_b_28,
	A_wr_data_unfiltered_2,
	A_wr_data_unfiltered_13,
	A_wr_data_unfiltered_12,
	A_wr_data_unfiltered_11,
	A_wr_data_unfiltered_10,
	A_wr_data_unfiltered_9,
	A_wr_data_unfiltered_8,
	A_wr_data_unfiltered_7,
	A_wr_data_unfiltered_6,
	A_wr_data_unfiltered_5,
	A_wr_data_unfiltered_4,
	A_wr_data_unfiltered_3,
	A_wr_data_unfiltered_1,
	A_wr_data_unfiltered_0,
	A_wr_data_unfiltered_21,
	A_wr_data_unfiltered_20,
	A_wr_data_unfiltered_25,
	A_wr_data_unfiltered_17,
	A_wr_data_unfiltered_24,
	A_wr_data_unfiltered_16,
	A_wr_data_unfiltered_27,
	A_wr_data_unfiltered_19,
	A_wr_data_unfiltered_26,
	A_wr_data_unfiltered_18,
	A_wr_data_unfiltered_23,
	A_wr_data_unfiltered_22,
	A_wr_data_unfiltered_29,
	A_wr_data_unfiltered_30,
	A_wr_data_unfiltered_31,
	A_wr_data_unfiltered_28,
	A_wr_data_unfiltered_15,
	A_wr_data_unfiltered_14,
	A_dst_regnum_from_M_4,
	A_wr_dst_reg_from_M,
	A_dst_regnum_from_M_0,
	A_dst_regnum_from_M_1,
	A_dst_regnum_from_M_2,
	A_dst_regnum_from_M_3,
	rf_b_rd_port_addr_0,
	rf_b_rd_port_addr_1,
	rf_b_rd_port_addr_2,
	rf_b_rd_port_addr_3,
	rf_b_rd_port_addr_4,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_b_2;
output 	q_b_13;
output 	q_b_12;
output 	q_b_11;
output 	q_b_10;
output 	q_b_9;
output 	q_b_8;
output 	q_b_7;
output 	q_b_6;
output 	q_b_5;
output 	q_b_4;
output 	q_b_3;
output 	q_b_1;
output 	q_b_0;
output 	q_b_21;
output 	q_b_20;
output 	q_b_25;
output 	q_b_17;
output 	q_b_24;
output 	q_b_16;
output 	q_b_27;
output 	q_b_19;
output 	q_b_26;
output 	q_b_18;
output 	q_b_23;
output 	q_b_15;
output 	q_b_22;
output 	q_b_14;
output 	q_b_29;
output 	q_b_30;
output 	q_b_31;
output 	q_b_28;
input 	A_wr_data_unfiltered_2;
input 	A_wr_data_unfiltered_13;
input 	A_wr_data_unfiltered_12;
input 	A_wr_data_unfiltered_11;
input 	A_wr_data_unfiltered_10;
input 	A_wr_data_unfiltered_9;
input 	A_wr_data_unfiltered_8;
input 	A_wr_data_unfiltered_7;
input 	A_wr_data_unfiltered_6;
input 	A_wr_data_unfiltered_5;
input 	A_wr_data_unfiltered_4;
input 	A_wr_data_unfiltered_3;
input 	A_wr_data_unfiltered_1;
input 	A_wr_data_unfiltered_0;
input 	A_wr_data_unfiltered_21;
input 	A_wr_data_unfiltered_20;
input 	A_wr_data_unfiltered_25;
input 	A_wr_data_unfiltered_17;
input 	A_wr_data_unfiltered_24;
input 	A_wr_data_unfiltered_16;
input 	A_wr_data_unfiltered_27;
input 	A_wr_data_unfiltered_19;
input 	A_wr_data_unfiltered_26;
input 	A_wr_data_unfiltered_18;
input 	A_wr_data_unfiltered_23;
input 	A_wr_data_unfiltered_22;
input 	A_wr_data_unfiltered_29;
input 	A_wr_data_unfiltered_30;
input 	A_wr_data_unfiltered_31;
input 	A_wr_data_unfiltered_28;
input 	A_wr_data_unfiltered_15;
input 	A_wr_data_unfiltered_14;
input 	A_dst_regnum_from_M_4;
input 	A_wr_dst_reg_from_M;
input 	A_dst_regnum_from_M_0;
input 	A_dst_regnum_from_M_1;
input 	A_dst_regnum_from_M_2;
input 	A_dst_regnum_from_M_3;
input 	rf_b_rd_port_addr_0;
input 	rf_b_rd_port_addr_1;
input 	rf_b_rd_port_addr_2;
input 	rf_b_rd_port_addr_3;
input 	rf_b_rd_port_addr_4;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_9 the_altsyncram(
	.q_b({q_b_31,q_b_30,q_b_29,q_b_28,q_b_27,q_b_26,q_b_25,q_b_24,q_b_23,q_b_22,q_b_21,q_b_20,q_b_19,q_b_18,q_b_17,q_b_16,q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.data_a({A_wr_data_unfiltered_31,A_wr_data_unfiltered_30,A_wr_data_unfiltered_29,A_wr_data_unfiltered_28,A_wr_data_unfiltered_27,A_wr_data_unfiltered_26,A_wr_data_unfiltered_25,A_wr_data_unfiltered_24,A_wr_data_unfiltered_23,A_wr_data_unfiltered_22,A_wr_data_unfiltered_21,
A_wr_data_unfiltered_20,A_wr_data_unfiltered_19,A_wr_data_unfiltered_18,A_wr_data_unfiltered_17,A_wr_data_unfiltered_16,A_wr_data_unfiltered_15,A_wr_data_unfiltered_14,A_wr_data_unfiltered_13,A_wr_data_unfiltered_12,A_wr_data_unfiltered_11,A_wr_data_unfiltered_10,
A_wr_data_unfiltered_9,A_wr_data_unfiltered_8,A_wr_data_unfiltered_7,A_wr_data_unfiltered_6,A_wr_data_unfiltered_5,A_wr_data_unfiltered_4,A_wr_data_unfiltered_3,A_wr_data_unfiltered_2,A_wr_data_unfiltered_1,A_wr_data_unfiltered_0}),
	.address_a({gnd,gnd,gnd,gnd,gnd,A_dst_regnum_from_M_4,A_dst_regnum_from_M_3,A_dst_regnum_from_M_2,A_dst_regnum_from_M_1,A_dst_regnum_from_M_0}),
	.wren_a(A_wr_dst_reg_from_M),
	.address_b({gnd,gnd,gnd,gnd,gnd,rf_b_rd_port_addr_4,rf_b_rd_port_addr_3,rf_b_rd_port_addr_2,rf_b_rd_port_addr_1,rf_b_rd_port_addr_0}),
	.clock0(clk_clk));

endmodule

module embedded_system_altsyncram_9 (
	q_b,
	data_a,
	address_a,
	wren_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	[9:0] address_a;
input 	wren_a;
input 	[9:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_atn1 auto_generated(
	.q_b({q_b[31],q_b[30],q_b[29],q_b[28],q_b[27],q_b[26],q_b[25],q_b[24],q_b[23],q_b[22],q_b[21],q_b[20],q_b[19],q_b[18],q_b[17],q_b[16],q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.wren_a(wren_a),
	.address_b({address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.clock0(clock0));

endmodule

module embedded_system_altsyncram_atn1 (
	q_b,
	data_a,
	address_a,
	wren_a,
	address_b,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_b;
input 	[31:0] data_a;
input 	[4:0] address_a;
input 	wren_a;
input 	[4:0] address_b;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a21_PORTBDATAOUT_bus;
wire [143:0] ram_block1a20_PORTBDATAOUT_bus;
wire [143:0] ram_block1a25_PORTBDATAOUT_bus;
wire [143:0] ram_block1a17_PORTBDATAOUT_bus;
wire [143:0] ram_block1a24_PORTBDATAOUT_bus;
wire [143:0] ram_block1a16_PORTBDATAOUT_bus;
wire [143:0] ram_block1a27_PORTBDATAOUT_bus;
wire [143:0] ram_block1a19_PORTBDATAOUT_bus;
wire [143:0] ram_block1a26_PORTBDATAOUT_bus;
wire [143:0] ram_block1a18_PORTBDATAOUT_bus;
wire [143:0] ram_block1a23_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a22_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a29_PORTBDATAOUT_bus;
wire [143:0] ram_block1a30_PORTBDATAOUT_bus;
wire [143:0] ram_block1a31_PORTBDATAOUT_bus;
wire [143:0] ram_block1a28_PORTBDATAOUT_bus;

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[21] = ram_block1a21_PORTBDATAOUT_bus[0];

assign q_b[20] = ram_block1a20_PORTBDATAOUT_bus[0];

assign q_b[25] = ram_block1a25_PORTBDATAOUT_bus[0];

assign q_b[17] = ram_block1a17_PORTBDATAOUT_bus[0];

assign q_b[24] = ram_block1a24_PORTBDATAOUT_bus[0];

assign q_b[16] = ram_block1a16_PORTBDATAOUT_bus[0];

assign q_b[27] = ram_block1a27_PORTBDATAOUT_bus[0];

assign q_b[19] = ram_block1a19_PORTBDATAOUT_bus[0];

assign q_b[26] = ram_block1a26_PORTBDATAOUT_bus[0];

assign q_b[18] = ram_block1a18_PORTBDATAOUT_bus[0];

assign q_b[23] = ram_block1a23_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[22] = ram_block1a22_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[29] = ram_block1a29_PORTBDATAOUT_bus[0];

assign q_b[30] = ram_block1a30_PORTBDATAOUT_bus[0];

assign q_b[31] = ram_block1a31_PORTBDATAOUT_bus[0];

assign q_b[28] = ram_block1a28_PORTBDATAOUT_bus[0];

cyclonev_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a2.init_file_layout = "port_b";
defparam ram_block1a2.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 5;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 31;
defparam ram_block1a2.port_a_logical_ram_depth = 32;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 5;
defparam ram_block1a2.port_b_data_out_clear = "none";
defparam ram_block1a2.port_b_data_out_clock = "none";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 31;
defparam ram_block1a2.port_b_logical_ram_depth = 32;
defparam ram_block1a2.port_b_logical_ram_width = 32;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a13.init_file_layout = "port_b";
defparam ram_block1a13.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 5;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 31;
defparam ram_block1a13.port_a_logical_ram_depth = 32;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_address_clear = "none";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 5;
defparam ram_block1a13.port_b_data_out_clear = "none";
defparam ram_block1a13.port_b_data_out_clock = "none";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 31;
defparam ram_block1a13.port_b_logical_ram_depth = 32;
defparam ram_block1a13.port_b_logical_ram_width = 32;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a12.init_file_layout = "port_b";
defparam ram_block1a12.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 5;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 31;
defparam ram_block1a12.port_a_logical_ram_depth = 32;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_address_clear = "none";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 5;
defparam ram_block1a12.port_b_data_out_clear = "none";
defparam ram_block1a12.port_b_data_out_clock = "none";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 31;
defparam ram_block1a12.port_b_logical_ram_depth = 32;
defparam ram_block1a12.port_b_logical_ram_width = 32;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a11.init_file_layout = "port_b";
defparam ram_block1a11.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 5;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 31;
defparam ram_block1a11.port_a_logical_ram_depth = 32;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_address_clear = "none";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 5;
defparam ram_block1a11.port_b_data_out_clear = "none";
defparam ram_block1a11.port_b_data_out_clock = "none";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 31;
defparam ram_block1a11.port_b_logical_ram_depth = 32;
defparam ram_block1a11.port_b_logical_ram_width = 32;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a10.init_file_layout = "port_b";
defparam ram_block1a10.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 5;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 31;
defparam ram_block1a10.port_a_logical_ram_depth = 32;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_address_clear = "none";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 5;
defparam ram_block1a10.port_b_data_out_clear = "none";
defparam ram_block1a10.port_b_data_out_clock = "none";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 31;
defparam ram_block1a10.port_b_logical_ram_depth = 32;
defparam ram_block1a10.port_b_logical_ram_width = 32;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a9.init_file_layout = "port_b";
defparam ram_block1a9.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 5;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 31;
defparam ram_block1a9.port_a_logical_ram_depth = 32;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_address_clear = "none";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 5;
defparam ram_block1a9.port_b_data_out_clear = "none";
defparam ram_block1a9.port_b_data_out_clock = "none";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 31;
defparam ram_block1a9.port_b_logical_ram_depth = 32;
defparam ram_block1a9.port_b_logical_ram_width = 32;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a8.init_file_layout = "port_b";
defparam ram_block1a8.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 5;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 31;
defparam ram_block1a8.port_a_logical_ram_depth = 32;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_address_clear = "none";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 5;
defparam ram_block1a8.port_b_data_out_clear = "none";
defparam ram_block1a8.port_b_data_out_clock = "none";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 31;
defparam ram_block1a8.port_b_logical_ram_depth = 32;
defparam ram_block1a8.port_b_logical_ram_width = 32;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a7.init_file_layout = "port_b";
defparam ram_block1a7.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 5;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 31;
defparam ram_block1a7.port_a_logical_ram_depth = 32;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 5;
defparam ram_block1a7.port_b_data_out_clear = "none";
defparam ram_block1a7.port_b_data_out_clock = "none";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 31;
defparam ram_block1a7.port_b_logical_ram_depth = 32;
defparam ram_block1a7.port_b_logical_ram_width = 32;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a6.init_file_layout = "port_b";
defparam ram_block1a6.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 5;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 31;
defparam ram_block1a6.port_a_logical_ram_depth = 32;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 5;
defparam ram_block1a6.port_b_data_out_clear = "none";
defparam ram_block1a6.port_b_data_out_clock = "none";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 31;
defparam ram_block1a6.port_b_logical_ram_depth = 32;
defparam ram_block1a6.port_b_logical_ram_width = 32;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a5.init_file_layout = "port_b";
defparam ram_block1a5.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 5;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 31;
defparam ram_block1a5.port_a_logical_ram_depth = 32;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 5;
defparam ram_block1a5.port_b_data_out_clear = "none";
defparam ram_block1a5.port_b_data_out_clock = "none";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 31;
defparam ram_block1a5.port_b_logical_ram_depth = 32;
defparam ram_block1a5.port_b_logical_ram_width = 32;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a4.init_file_layout = "port_b";
defparam ram_block1a4.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 5;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 31;
defparam ram_block1a4.port_a_logical_ram_depth = 32;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 5;
defparam ram_block1a4.port_b_data_out_clear = "none";
defparam ram_block1a4.port_b_data_out_clock = "none";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 31;
defparam ram_block1a4.port_b_logical_ram_depth = 32;
defparam ram_block1a4.port_b_logical_ram_width = 32;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a3.init_file_layout = "port_b";
defparam ram_block1a3.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 5;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 31;
defparam ram_block1a3.port_a_logical_ram_depth = 32;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 5;
defparam ram_block1a3.port_b_data_out_clear = "none";
defparam ram_block1a3.port_b_data_out_clock = "none";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 31;
defparam ram_block1a3.port_b_logical_ram_depth = 32;
defparam ram_block1a3.port_b_logical_ram_width = 32;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a1.init_file_layout = "port_b";
defparam ram_block1a1.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 5;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 31;
defparam ram_block1a1.port_a_logical_ram_depth = 32;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 5;
defparam ram_block1a1.port_b_data_out_clear = "none";
defparam ram_block1a1.port_b_data_out_clock = "none";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 31;
defparam ram_block1a1.port_b_logical_ram_depth = 32;
defparam ram_block1a1.port_b_logical_ram_width = 32;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a0.init_file_layout = "port_b";
defparam ram_block1a0.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 5;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 31;
defparam ram_block1a0.port_a_logical_ram_depth = 32;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 5;
defparam ram_block1a0.port_b_data_out_clear = "none";
defparam ram_block1a0.port_b_data_out_clock = "none";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 31;
defparam ram_block1a0.port_b_logical_ram_depth = 32;
defparam ram_block1a0.port_b_logical_ram_width = 32;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a21(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a21_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a21.init_file_layout = "port_b";
defparam ram_block1a21.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.mixed_port_feed_through_mode = "old";
defparam ram_block1a21.operation_mode = "dual_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 5;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 31;
defparam ram_block1a21.port_a_logical_ram_depth = 32;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_address_clear = "none";
defparam ram_block1a21.port_b_address_clock = "clock0";
defparam ram_block1a21.port_b_address_width = 5;
defparam ram_block1a21.port_b_data_out_clear = "none";
defparam ram_block1a21.port_b_data_out_clock = "none";
defparam ram_block1a21.port_b_data_width = 1;
defparam ram_block1a21.port_b_first_address = 0;
defparam ram_block1a21.port_b_first_bit_number = 21;
defparam ram_block1a21.port_b_last_address = 31;
defparam ram_block1a21.port_b_logical_ram_depth = 32;
defparam ram_block1a21.port_b_logical_ram_width = 32;
defparam ram_block1a21.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a21.port_b_read_enable_clock = "clock0";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a20(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a20_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a20.init_file_layout = "port_b";
defparam ram_block1a20.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.mixed_port_feed_through_mode = "old";
defparam ram_block1a20.operation_mode = "dual_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 5;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 31;
defparam ram_block1a20.port_a_logical_ram_depth = 32;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_address_clear = "none";
defparam ram_block1a20.port_b_address_clock = "clock0";
defparam ram_block1a20.port_b_address_width = 5;
defparam ram_block1a20.port_b_data_out_clear = "none";
defparam ram_block1a20.port_b_data_out_clock = "none";
defparam ram_block1a20.port_b_data_width = 1;
defparam ram_block1a20.port_b_first_address = 0;
defparam ram_block1a20.port_b_first_bit_number = 20;
defparam ram_block1a20.port_b_last_address = 31;
defparam ram_block1a20.port_b_logical_ram_depth = 32;
defparam ram_block1a20.port_b_logical_ram_width = 32;
defparam ram_block1a20.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a20.port_b_read_enable_clock = "clock0";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a25(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a25_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a25.init_file_layout = "port_b";
defparam ram_block1a25.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.mixed_port_feed_through_mode = "old";
defparam ram_block1a25.operation_mode = "dual_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 5;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 31;
defparam ram_block1a25.port_a_logical_ram_depth = 32;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_address_clear = "none";
defparam ram_block1a25.port_b_address_clock = "clock0";
defparam ram_block1a25.port_b_address_width = 5;
defparam ram_block1a25.port_b_data_out_clear = "none";
defparam ram_block1a25.port_b_data_out_clock = "none";
defparam ram_block1a25.port_b_data_width = 1;
defparam ram_block1a25.port_b_first_address = 0;
defparam ram_block1a25.port_b_first_bit_number = 25;
defparam ram_block1a25.port_b_last_address = 31;
defparam ram_block1a25.port_b_logical_ram_depth = 32;
defparam ram_block1a25.port_b_logical_ram_width = 32;
defparam ram_block1a25.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a25.port_b_read_enable_clock = "clock0";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a17(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a17_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a17.init_file_layout = "port_b";
defparam ram_block1a17.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.mixed_port_feed_through_mode = "old";
defparam ram_block1a17.operation_mode = "dual_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 5;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 31;
defparam ram_block1a17.port_a_logical_ram_depth = 32;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_address_clear = "none";
defparam ram_block1a17.port_b_address_clock = "clock0";
defparam ram_block1a17.port_b_address_width = 5;
defparam ram_block1a17.port_b_data_out_clear = "none";
defparam ram_block1a17.port_b_data_out_clock = "none";
defparam ram_block1a17.port_b_data_width = 1;
defparam ram_block1a17.port_b_first_address = 0;
defparam ram_block1a17.port_b_first_bit_number = 17;
defparam ram_block1a17.port_b_last_address = 31;
defparam ram_block1a17.port_b_logical_ram_depth = 32;
defparam ram_block1a17.port_b_logical_ram_width = 32;
defparam ram_block1a17.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a17.port_b_read_enable_clock = "clock0";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a24(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a24_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a24.init_file_layout = "port_b";
defparam ram_block1a24.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.mixed_port_feed_through_mode = "old";
defparam ram_block1a24.operation_mode = "dual_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 5;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 31;
defparam ram_block1a24.port_a_logical_ram_depth = 32;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_address_clear = "none";
defparam ram_block1a24.port_b_address_clock = "clock0";
defparam ram_block1a24.port_b_address_width = 5;
defparam ram_block1a24.port_b_data_out_clear = "none";
defparam ram_block1a24.port_b_data_out_clock = "none";
defparam ram_block1a24.port_b_data_width = 1;
defparam ram_block1a24.port_b_first_address = 0;
defparam ram_block1a24.port_b_first_bit_number = 24;
defparam ram_block1a24.port_b_last_address = 31;
defparam ram_block1a24.port_b_logical_ram_depth = 32;
defparam ram_block1a24.port_b_logical_ram_width = 32;
defparam ram_block1a24.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a24.port_b_read_enable_clock = "clock0";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a16(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a16_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a16.init_file_layout = "port_b";
defparam ram_block1a16.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.mixed_port_feed_through_mode = "old";
defparam ram_block1a16.operation_mode = "dual_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 5;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 31;
defparam ram_block1a16.port_a_logical_ram_depth = 32;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_address_clear = "none";
defparam ram_block1a16.port_b_address_clock = "clock0";
defparam ram_block1a16.port_b_address_width = 5;
defparam ram_block1a16.port_b_data_out_clear = "none";
defparam ram_block1a16.port_b_data_out_clock = "none";
defparam ram_block1a16.port_b_data_width = 1;
defparam ram_block1a16.port_b_first_address = 0;
defparam ram_block1a16.port_b_first_bit_number = 16;
defparam ram_block1a16.port_b_last_address = 31;
defparam ram_block1a16.port_b_logical_ram_depth = 32;
defparam ram_block1a16.port_b_logical_ram_width = 32;
defparam ram_block1a16.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a16.port_b_read_enable_clock = "clock0";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a27(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a27_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a27.init_file_layout = "port_b";
defparam ram_block1a27.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.mixed_port_feed_through_mode = "old";
defparam ram_block1a27.operation_mode = "dual_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 5;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 31;
defparam ram_block1a27.port_a_logical_ram_depth = 32;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_address_clear = "none";
defparam ram_block1a27.port_b_address_clock = "clock0";
defparam ram_block1a27.port_b_address_width = 5;
defparam ram_block1a27.port_b_data_out_clear = "none";
defparam ram_block1a27.port_b_data_out_clock = "none";
defparam ram_block1a27.port_b_data_width = 1;
defparam ram_block1a27.port_b_first_address = 0;
defparam ram_block1a27.port_b_first_bit_number = 27;
defparam ram_block1a27.port_b_last_address = 31;
defparam ram_block1a27.port_b_logical_ram_depth = 32;
defparam ram_block1a27.port_b_logical_ram_width = 32;
defparam ram_block1a27.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a27.port_b_read_enable_clock = "clock0";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a19(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a19_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a19.init_file_layout = "port_b";
defparam ram_block1a19.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.mixed_port_feed_through_mode = "old";
defparam ram_block1a19.operation_mode = "dual_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 5;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 31;
defparam ram_block1a19.port_a_logical_ram_depth = 32;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_address_clear = "none";
defparam ram_block1a19.port_b_address_clock = "clock0";
defparam ram_block1a19.port_b_address_width = 5;
defparam ram_block1a19.port_b_data_out_clear = "none";
defparam ram_block1a19.port_b_data_out_clock = "none";
defparam ram_block1a19.port_b_data_width = 1;
defparam ram_block1a19.port_b_first_address = 0;
defparam ram_block1a19.port_b_first_bit_number = 19;
defparam ram_block1a19.port_b_last_address = 31;
defparam ram_block1a19.port_b_logical_ram_depth = 32;
defparam ram_block1a19.port_b_logical_ram_width = 32;
defparam ram_block1a19.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a19.port_b_read_enable_clock = "clock0";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a26(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a26_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a26.init_file_layout = "port_b";
defparam ram_block1a26.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.mixed_port_feed_through_mode = "old";
defparam ram_block1a26.operation_mode = "dual_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 5;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 31;
defparam ram_block1a26.port_a_logical_ram_depth = 32;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_address_clear = "none";
defparam ram_block1a26.port_b_address_clock = "clock0";
defparam ram_block1a26.port_b_address_width = 5;
defparam ram_block1a26.port_b_data_out_clear = "none";
defparam ram_block1a26.port_b_data_out_clock = "none";
defparam ram_block1a26.port_b_data_width = 1;
defparam ram_block1a26.port_b_first_address = 0;
defparam ram_block1a26.port_b_first_bit_number = 26;
defparam ram_block1a26.port_b_last_address = 31;
defparam ram_block1a26.port_b_logical_ram_depth = 32;
defparam ram_block1a26.port_b_logical_ram_width = 32;
defparam ram_block1a26.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a26.port_b_read_enable_clock = "clock0";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a18(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a18_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a18.init_file_layout = "port_b";
defparam ram_block1a18.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.mixed_port_feed_through_mode = "old";
defparam ram_block1a18.operation_mode = "dual_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 5;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 31;
defparam ram_block1a18.port_a_logical_ram_depth = 32;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_address_clear = "none";
defparam ram_block1a18.port_b_address_clock = "clock0";
defparam ram_block1a18.port_b_address_width = 5;
defparam ram_block1a18.port_b_data_out_clear = "none";
defparam ram_block1a18.port_b_data_out_clock = "none";
defparam ram_block1a18.port_b_data_width = 1;
defparam ram_block1a18.port_b_first_address = 0;
defparam ram_block1a18.port_b_first_bit_number = 18;
defparam ram_block1a18.port_b_last_address = 31;
defparam ram_block1a18.port_b_logical_ram_depth = 32;
defparam ram_block1a18.port_b_logical_ram_width = 32;
defparam ram_block1a18.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a18.port_b_read_enable_clock = "clock0";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a23(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a23_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a23.init_file_layout = "port_b";
defparam ram_block1a23.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.mixed_port_feed_through_mode = "old";
defparam ram_block1a23.operation_mode = "dual_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 5;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 31;
defparam ram_block1a23.port_a_logical_ram_depth = 32;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_address_clear = "none";
defparam ram_block1a23.port_b_address_clock = "clock0";
defparam ram_block1a23.port_b_address_width = 5;
defparam ram_block1a23.port_b_data_out_clear = "none";
defparam ram_block1a23.port_b_data_out_clock = "none";
defparam ram_block1a23.port_b_data_width = 1;
defparam ram_block1a23.port_b_first_address = 0;
defparam ram_block1a23.port_b_first_bit_number = 23;
defparam ram_block1a23.port_b_last_address = 31;
defparam ram_block1a23.port_b_logical_ram_depth = 32;
defparam ram_block1a23.port_b_logical_ram_width = 32;
defparam ram_block1a23.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a23.port_b_read_enable_clock = "clock0";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a15.init_file_layout = "port_b";
defparam ram_block1a15.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 5;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 31;
defparam ram_block1a15.port_a_logical_ram_depth = 32;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_address_clear = "none";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 5;
defparam ram_block1a15.port_b_data_out_clear = "none";
defparam ram_block1a15.port_b_data_out_clock = "none";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 31;
defparam ram_block1a15.port_b_logical_ram_depth = 32;
defparam ram_block1a15.port_b_logical_ram_width = 32;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a22(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a22_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a22.init_file_layout = "port_b";
defparam ram_block1a22.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.mixed_port_feed_through_mode = "old";
defparam ram_block1a22.operation_mode = "dual_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 5;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 31;
defparam ram_block1a22.port_a_logical_ram_depth = 32;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_address_clear = "none";
defparam ram_block1a22.port_b_address_clock = "clock0";
defparam ram_block1a22.port_b_address_width = 5;
defparam ram_block1a22.port_b_data_out_clear = "none";
defparam ram_block1a22.port_b_data_out_clock = "none";
defparam ram_block1a22.port_b_data_width = 1;
defparam ram_block1a22.port_b_first_address = 0;
defparam ram_block1a22.port_b_first_bit_number = 22;
defparam ram_block1a22.port_b_last_address = 31;
defparam ram_block1a22.port_b_logical_ram_depth = 32;
defparam ram_block1a22.port_b_logical_ram_width = 32;
defparam ram_block1a22.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a22.port_b_read_enable_clock = "clock0";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a14.init_file_layout = "port_b";
defparam ram_block1a14.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 5;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 31;
defparam ram_block1a14.port_a_logical_ram_depth = 32;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_address_clear = "none";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 5;
defparam ram_block1a14.port_b_data_out_clear = "none";
defparam ram_block1a14.port_b_data_out_clock = "none";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 31;
defparam ram_block1a14.port_b_logical_ram_depth = 32;
defparam ram_block1a14.port_b_logical_ram_width = 32;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a29(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a29_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a29.init_file_layout = "port_b";
defparam ram_block1a29.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.mixed_port_feed_through_mode = "old";
defparam ram_block1a29.operation_mode = "dual_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 5;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 31;
defparam ram_block1a29.port_a_logical_ram_depth = 32;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_address_clear = "none";
defparam ram_block1a29.port_b_address_clock = "clock0";
defparam ram_block1a29.port_b_address_width = 5;
defparam ram_block1a29.port_b_data_out_clear = "none";
defparam ram_block1a29.port_b_data_out_clock = "none";
defparam ram_block1a29.port_b_data_width = 1;
defparam ram_block1a29.port_b_first_address = 0;
defparam ram_block1a29.port_b_first_bit_number = 29;
defparam ram_block1a29.port_b_last_address = 31;
defparam ram_block1a29.port_b_logical_ram_depth = 32;
defparam ram_block1a29.port_b_logical_ram_width = 32;
defparam ram_block1a29.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a29.port_b_read_enable_clock = "clock0";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = "00000000";

cyclonev_ram_block ram_block1a30(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a30_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a30.init_file_layout = "port_b";
defparam ram_block1a30.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.mixed_port_feed_through_mode = "old";
defparam ram_block1a30.operation_mode = "dual_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 5;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 31;
defparam ram_block1a30.port_a_logical_ram_depth = 32;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_address_clear = "none";
defparam ram_block1a30.port_b_address_clock = "clock0";
defparam ram_block1a30.port_b_address_width = 5;
defparam ram_block1a30.port_b_data_out_clear = "none";
defparam ram_block1a30.port_b_data_out_clock = "none";
defparam ram_block1a30.port_b_data_width = 1;
defparam ram_block1a30.port_b_first_address = 0;
defparam ram_block1a30.port_b_first_bit_number = 30;
defparam ram_block1a30.port_b_last_address = 31;
defparam ram_block1a30.port_b_logical_ram_depth = 32;
defparam ram_block1a30.port_b_logical_ram_width = 32;
defparam ram_block1a30.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a30.port_b_read_enable_clock = "clock0";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a31(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a31_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a31.init_file_layout = "port_b";
defparam ram_block1a31.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.mixed_port_feed_through_mode = "old";
defparam ram_block1a31.operation_mode = "dual_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 5;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 31;
defparam ram_block1a31.port_a_logical_ram_depth = 32;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_address_clear = "none";
defparam ram_block1a31.port_b_address_clock = "clock0";
defparam ram_block1a31.port_b_address_width = 5;
defparam ram_block1a31.port_b_data_out_clear = "none";
defparam ram_block1a31.port_b_data_out_clock = "none";
defparam ram_block1a31.port_b_data_width = 1;
defparam ram_block1a31.port_b_first_address = 0;
defparam ram_block1a31.port_b_first_bit_number = 31;
defparam ram_block1a31.port_b_last_address = 31;
defparam ram_block1a31.port_b_logical_ram_depth = 32;
defparam ram_block1a31.port_b_logical_ram_width = 32;
defparam ram_block1a31.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a31.port_b_read_enable_clock = "clock0";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = "FFFFFFFF";

cyclonev_ram_block ram_block1a28(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(vcc),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a28_PORTBDATAOUT_bus),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "embedded_system_nios2_qsys_0_rf_ram_b.mif";
defparam ram_block1a28.init_file_layout = "port_b";
defparam ram_block1a28.logical_ram_name = "embedded_system_nios2_qsys_0:nios2_qsys_0|embedded_system_nios2_qsys_0_register_bank_b_module:embedded_system_nios2_qsys_0_register_bank_b|altsyncram:the_altsyncram|altsyncram_atn1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.mixed_port_feed_through_mode = "old";
defparam ram_block1a28.operation_mode = "dual_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 5;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 31;
defparam ram_block1a28.port_a_logical_ram_depth = 32;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_address_clear = "none";
defparam ram_block1a28.port_b_address_clock = "clock0";
defparam ram_block1a28.port_b_address_width = 5;
defparam ram_block1a28.port_b_data_out_clear = "none";
defparam ram_block1a28.port_b_data_out_clock = "none";
defparam ram_block1a28.port_b_data_width = 1;
defparam ram_block1a28.port_b_first_address = 0;
defparam ram_block1a28.port_b_first_bit_number = 28;
defparam ram_block1a28.port_b_last_address = 31;
defparam ram_block1a28.port_b_logical_ram_depth = 32;
defparam ram_block1a28.port_b_logical_ram_width = 32;
defparam ram_block1a28.port_b_read_during_write_mode = "new_data_no_nbe_read";
defparam ram_block1a28.port_b_read_enable_clock = "clock0";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = "FFFFFFFF";

endmodule

module embedded_system_embedded_system_onchip_memory2_0 (
	q_a_2,
	q_a_10,
	q_a_18,
	q_a_26,
	q_a_7,
	q_a_23,
	q_a_15,
	q_a_31,
	q_a_29,
	q_a_13,
	q_a_28,
	q_a_12,
	q_a_27,
	q_a_11,
	q_a_25,
	q_a_9,
	q_a_24,
	q_a_8,
	q_a_6,
	q_a_14,
	q_a_22,
	q_a_30,
	q_a_5,
	q_a_21,
	q_a_4,
	q_a_20,
	q_a_3,
	q_a_19,
	q_a_1,
	q_a_17,
	q_a_0,
	q_a_16,
	d_write,
	saved_grant_0,
	mem_used_1,
	src1_valid,
	src2_valid,
	saved_grant_1,
	r_early_rst,
	src_payload,
	src_data_38,
	src_data_39,
	src_data_40,
	src_data_41,
	src_data_42,
	src_data_43,
	src_data_44,
	src_data_45,
	src_data_46,
	src_data_47,
	src_data_32,
	src_payload1,
	src_data_33,
	src_payload2,
	src_data_34,
	src_payload3,
	src_data_35,
	src_payload4,
	src_payload5,
	src_payload6,
	src_payload7,
	src_payload8,
	src_payload9,
	src_payload10,
	src_payload11,
	src_payload12,
	src_payload13,
	src_payload14,
	src_payload15,
	src_payload16,
	src_payload17,
	src_payload18,
	src_payload19,
	src_payload20,
	src_payload21,
	src_payload22,
	src_payload23,
	src_payload24,
	src_payload25,
	src_payload26,
	src_payload27,
	src_payload28,
	src_payload29,
	src_payload30,
	src_payload31,
	clk_clk)/* synthesis synthesis_greybox=1 */;
output 	q_a_2;
output 	q_a_10;
output 	q_a_18;
output 	q_a_26;
output 	q_a_7;
output 	q_a_23;
output 	q_a_15;
output 	q_a_31;
output 	q_a_29;
output 	q_a_13;
output 	q_a_28;
output 	q_a_12;
output 	q_a_27;
output 	q_a_11;
output 	q_a_25;
output 	q_a_9;
output 	q_a_24;
output 	q_a_8;
output 	q_a_6;
output 	q_a_14;
output 	q_a_22;
output 	q_a_30;
output 	q_a_5;
output 	q_a_21;
output 	q_a_4;
output 	q_a_20;
output 	q_a_3;
output 	q_a_19;
output 	q_a_1;
output 	q_a_17;
output 	q_a_0;
output 	q_a_16;
input 	d_write;
input 	saved_grant_0;
input 	mem_used_1;
input 	src1_valid;
input 	src2_valid;
input 	saved_grant_1;
input 	r_early_rst;
input 	src_payload;
input 	src_data_38;
input 	src_data_39;
input 	src_data_40;
input 	src_data_41;
input 	src_data_42;
input 	src_data_43;
input 	src_data_44;
input 	src_data_45;
input 	src_data_46;
input 	src_data_47;
input 	src_data_32;
input 	src_payload1;
input 	src_data_33;
input 	src_payload2;
input 	src_data_34;
input 	src_payload3;
input 	src_data_35;
input 	src_payload4;
input 	src_payload5;
input 	src_payload6;
input 	src_payload7;
input 	src_payload8;
input 	src_payload9;
input 	src_payload10;
input 	src_payload11;
input 	src_payload12;
input 	src_payload13;
input 	src_payload14;
input 	src_payload15;
input 	src_payload16;
input 	src_payload17;
input 	src_payload18;
input 	src_payload19;
input 	src_payload20;
input 	src_payload21;
input 	src_payload22;
input 	src_payload23;
input 	src_payload24;
input 	src_payload25;
input 	src_payload26;
input 	src_payload27;
input 	src_payload28;
input 	src_payload29;
input 	src_payload30;
input 	src_payload31;
input 	clk_clk;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wren~0_combout ;


embedded_system_altsyncram_10 the_altsyncram(
	.q_a({q_a_31,q_a_30,q_a_29,q_a_28,q_a_27,q_a_26,q_a_25,q_a_24,q_a_23,q_a_22,q_a_21,q_a_20,q_a_19,q_a_18,q_a_17,q_a_16,q_a_15,q_a_14,q_a_13,q_a_12,q_a_11,q_a_10,q_a_9,q_a_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.clocken0(r_early_rst),
	.wren_a(\wren~0_combout ),
	.data_a({src_payload7,src_payload21,src_payload8,src_payload10,src_payload12,src_payload3,src_payload14,src_payload16,src_payload5,src_payload20,src_payload23,src_payload25,src_payload27,src_payload2,src_payload29,src_payload31,src_payload6,src_payload19,src_payload9,src_payload11,
src_payload13,src_payload1,src_payload15,src_payload17,src_payload4,src_payload18,src_payload22,src_payload24,src_payload26,src_payload,src_payload28,src_payload30}),
	.address_a({src_data_47,src_data_46,src_data_45,src_data_44,src_data_43,src_data_42,src_data_41,src_data_40,src_data_39,src_data_38}),
	.byteena_a({src_data_35,src_data_34,src_data_33,src_data_32}),
	.clock0(clk_clk));

cyclonev_lcell_comb \wren~0 (
	.dataa(!d_write),
	.datab(!saved_grant_0),
	.datac(!mem_used_1),
	.datad(!src1_valid),
	.datae(!src2_valid),
	.dataf(!saved_grant_1),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\wren~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \wren~0 .extended_lut = "off";
defparam \wren~0 .lut_mask = 64'hFFFFFFFFFFFFFFEF;
defparam \wren~0 .shared_arith = "off";

endmodule

module embedded_system_altsyncram_10 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[9:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



embedded_system_altsyncram_45o1 auto_generated(
	.q_a({q_a[31],q_a[30],q_a[29],q_a[28],q_a[27],q_a[26],q_a[25],q_a[24],q_a[23],q_a[22],q_a[21],q_a[20],q_a[19],q_a[18],q_a[17],q_a[16],q_a[15],q_a[14],q_a[13],q_a[12],q_a[11],q_a[10],q_a[9],q_a[8],q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.clocken0(clocken0),
	.wren_a(wren_a),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_a({address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.byteena_a({byteena_a[3],byteena_a[2],byteena_a[1],byteena_a[0]}),
	.clock0(clock0));

endmodule

module embedded_system_altsyncram_45o1 (
	q_a,
	clocken0,
	wren_a,
	data_a,
	address_a,
	byteena_a,
	clock0)/* synthesis synthesis_greybox=1 */;
output 	[31:0] q_a;
input 	clocken0;
input 	wren_a;
input 	[31:0] data_a;
input 	[9:0] address_a;
input 	[3:0] byteena_a;
input 	clock0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a10_PORTADATAOUT_bus;
wire [143:0] ram_block1a18_PORTADATAOUT_bus;
wire [143:0] ram_block1a26_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a23_PORTADATAOUT_bus;
wire [143:0] ram_block1a15_PORTADATAOUT_bus;
wire [143:0] ram_block1a31_PORTADATAOUT_bus;
wire [143:0] ram_block1a29_PORTADATAOUT_bus;
wire [143:0] ram_block1a13_PORTADATAOUT_bus;
wire [143:0] ram_block1a28_PORTADATAOUT_bus;
wire [143:0] ram_block1a12_PORTADATAOUT_bus;
wire [143:0] ram_block1a27_PORTADATAOUT_bus;
wire [143:0] ram_block1a11_PORTADATAOUT_bus;
wire [143:0] ram_block1a25_PORTADATAOUT_bus;
wire [143:0] ram_block1a9_PORTADATAOUT_bus;
wire [143:0] ram_block1a24_PORTADATAOUT_bus;
wire [143:0] ram_block1a8_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a14_PORTADATAOUT_bus;
wire [143:0] ram_block1a22_PORTADATAOUT_bus;
wire [143:0] ram_block1a30_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a21_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a20_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a19_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a17_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a16_PORTADATAOUT_bus;

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_a[10] = ram_block1a10_PORTADATAOUT_bus[0];

assign q_a[18] = ram_block1a18_PORTADATAOUT_bus[0];

assign q_a[26] = ram_block1a26_PORTADATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_a[23] = ram_block1a23_PORTADATAOUT_bus[0];

assign q_a[15] = ram_block1a15_PORTADATAOUT_bus[0];

assign q_a[31] = ram_block1a31_PORTADATAOUT_bus[0];

assign q_a[29] = ram_block1a29_PORTADATAOUT_bus[0];

assign q_a[13] = ram_block1a13_PORTADATAOUT_bus[0];

assign q_a[28] = ram_block1a28_PORTADATAOUT_bus[0];

assign q_a[12] = ram_block1a12_PORTADATAOUT_bus[0];

assign q_a[27] = ram_block1a27_PORTADATAOUT_bus[0];

assign q_a[11] = ram_block1a11_PORTADATAOUT_bus[0];

assign q_a[25] = ram_block1a25_PORTADATAOUT_bus[0];

assign q_a[9] = ram_block1a9_PORTADATAOUT_bus[0];

assign q_a[24] = ram_block1a24_PORTADATAOUT_bus[0];

assign q_a[8] = ram_block1a8_PORTADATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_a[14] = ram_block1a14_PORTADATAOUT_bus[0];

assign q_a[22] = ram_block1a22_PORTADATAOUT_bus[0];

assign q_a[30] = ram_block1a30_PORTADATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_a[21] = ram_block1a21_PORTADATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_a[20] = ram_block1a20_PORTADATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_a[19] = ram_block1a19_PORTADATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_a[17] = ram_block1a17_PORTADATAOUT_bus[0];

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_a[16] = ram_block1a16_PORTADATAOUT_bus[0];

cyclonev_ram_block ram_block1a2(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.operation_mode = "single_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 10;
defparam ram_block1a2.port_a_byte_enable_mask_width = 1;
defparam ram_block1a2.port_a_byte_size = 1;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 1023;
defparam ram_block1a2.port_a_logical_ram_depth = 1024;
defparam ram_block1a2.port_a_logical_ram_width = 32;
defparam ram_block1a2.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a10(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a10_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a10.init_file_layout = "port_a";
defparam ram_block1a10.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.operation_mode = "single_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 10;
defparam ram_block1a10.port_a_byte_enable_mask_width = 1;
defparam ram_block1a10.port_a_byte_size = 1;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 1023;
defparam ram_block1a10.port_a_logical_ram_depth = 1024;
defparam ram_block1a10.port_a_logical_ram_width = 32;
defparam ram_block1a10.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a10.ram_block_type = "auto";
defparam ram_block1a10.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a18(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[18]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a18_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a18.clk0_core_clock_enable = "ena0";
defparam ram_block1a18.clk0_input_clock_enable = "ena0";
defparam ram_block1a18.data_interleave_offset_in_bits = 1;
defparam ram_block1a18.data_interleave_width_in_bits = 1;
defparam ram_block1a18.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a18.init_file_layout = "port_a";
defparam ram_block1a18.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a18.operation_mode = "single_port";
defparam ram_block1a18.port_a_address_clear = "none";
defparam ram_block1a18.port_a_address_width = 10;
defparam ram_block1a18.port_a_byte_enable_mask_width = 1;
defparam ram_block1a18.port_a_byte_size = 1;
defparam ram_block1a18.port_a_data_out_clear = "none";
defparam ram_block1a18.port_a_data_out_clock = "none";
defparam ram_block1a18.port_a_data_width = 1;
defparam ram_block1a18.port_a_first_address = 0;
defparam ram_block1a18.port_a_first_bit_number = 18;
defparam ram_block1a18.port_a_last_address = 1023;
defparam ram_block1a18.port_a_logical_ram_depth = 1024;
defparam ram_block1a18.port_a_logical_ram_width = 32;
defparam ram_block1a18.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a18.ram_block_type = "auto";
defparam ram_block1a18.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a26(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[26]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a26_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a26.clk0_core_clock_enable = "ena0";
defparam ram_block1a26.clk0_input_clock_enable = "ena0";
defparam ram_block1a26.data_interleave_offset_in_bits = 1;
defparam ram_block1a26.data_interleave_width_in_bits = 1;
defparam ram_block1a26.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a26.init_file_layout = "port_a";
defparam ram_block1a26.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a26.operation_mode = "single_port";
defparam ram_block1a26.port_a_address_clear = "none";
defparam ram_block1a26.port_a_address_width = 10;
defparam ram_block1a26.port_a_byte_enable_mask_width = 1;
defparam ram_block1a26.port_a_byte_size = 1;
defparam ram_block1a26.port_a_data_out_clear = "none";
defparam ram_block1a26.port_a_data_out_clock = "none";
defparam ram_block1a26.port_a_data_width = 1;
defparam ram_block1a26.port_a_first_address = 0;
defparam ram_block1a26.port_a_first_bit_number = 26;
defparam ram_block1a26.port_a_last_address = 1023;
defparam ram_block1a26.port_a_logical_ram_depth = 1024;
defparam ram_block1a26.port_a_logical_ram_width = 32;
defparam ram_block1a26.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a26.ram_block_type = "auto";
defparam ram_block1a26.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a7(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.operation_mode = "single_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 10;
defparam ram_block1a7.port_a_byte_enable_mask_width = 1;
defparam ram_block1a7.port_a_byte_size = 1;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 1023;
defparam ram_block1a7.port_a_logical_ram_depth = 1024;
defparam ram_block1a7.port_a_logical_ram_width = 32;
defparam ram_block1a7.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a23(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[23]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a23_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a23.clk0_core_clock_enable = "ena0";
defparam ram_block1a23.clk0_input_clock_enable = "ena0";
defparam ram_block1a23.data_interleave_offset_in_bits = 1;
defparam ram_block1a23.data_interleave_width_in_bits = 1;
defparam ram_block1a23.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a23.init_file_layout = "port_a";
defparam ram_block1a23.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a23.operation_mode = "single_port";
defparam ram_block1a23.port_a_address_clear = "none";
defparam ram_block1a23.port_a_address_width = 10;
defparam ram_block1a23.port_a_byte_enable_mask_width = 1;
defparam ram_block1a23.port_a_byte_size = 1;
defparam ram_block1a23.port_a_data_out_clear = "none";
defparam ram_block1a23.port_a_data_out_clock = "none";
defparam ram_block1a23.port_a_data_width = 1;
defparam ram_block1a23.port_a_first_address = 0;
defparam ram_block1a23.port_a_first_bit_number = 23;
defparam ram_block1a23.port_a_last_address = 1023;
defparam ram_block1a23.port_a_logical_ram_depth = 1024;
defparam ram_block1a23.port_a_logical_ram_width = 32;
defparam ram_block1a23.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a23.ram_block_type = "auto";
defparam ram_block1a23.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a15(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a15_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a15.init_file_layout = "port_a";
defparam ram_block1a15.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.operation_mode = "single_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 10;
defparam ram_block1a15.port_a_byte_enable_mask_width = 1;
defparam ram_block1a15.port_a_byte_size = 1;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 1023;
defparam ram_block1a15.port_a_logical_ram_depth = 1024;
defparam ram_block1a15.port_a_logical_ram_width = 32;
defparam ram_block1a15.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a15.ram_block_type = "auto";
defparam ram_block1a15.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a31(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[31]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a31_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a31.clk0_core_clock_enable = "ena0";
defparam ram_block1a31.clk0_input_clock_enable = "ena0";
defparam ram_block1a31.data_interleave_offset_in_bits = 1;
defparam ram_block1a31.data_interleave_width_in_bits = 1;
defparam ram_block1a31.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a31.init_file_layout = "port_a";
defparam ram_block1a31.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a31.operation_mode = "single_port";
defparam ram_block1a31.port_a_address_clear = "none";
defparam ram_block1a31.port_a_address_width = 10;
defparam ram_block1a31.port_a_byte_enable_mask_width = 1;
defparam ram_block1a31.port_a_byte_size = 1;
defparam ram_block1a31.port_a_data_out_clear = "none";
defparam ram_block1a31.port_a_data_out_clock = "none";
defparam ram_block1a31.port_a_data_width = 1;
defparam ram_block1a31.port_a_first_address = 0;
defparam ram_block1a31.port_a_first_bit_number = 31;
defparam ram_block1a31.port_a_last_address = 1023;
defparam ram_block1a31.port_a_logical_ram_depth = 1024;
defparam ram_block1a31.port_a_logical_ram_width = 32;
defparam ram_block1a31.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a31.ram_block_type = "auto";
defparam ram_block1a31.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a29(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[29]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a29_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a29.clk0_core_clock_enable = "ena0";
defparam ram_block1a29.clk0_input_clock_enable = "ena0";
defparam ram_block1a29.data_interleave_offset_in_bits = 1;
defparam ram_block1a29.data_interleave_width_in_bits = 1;
defparam ram_block1a29.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a29.init_file_layout = "port_a";
defparam ram_block1a29.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a29.operation_mode = "single_port";
defparam ram_block1a29.port_a_address_clear = "none";
defparam ram_block1a29.port_a_address_width = 10;
defparam ram_block1a29.port_a_byte_enable_mask_width = 1;
defparam ram_block1a29.port_a_byte_size = 1;
defparam ram_block1a29.port_a_data_out_clear = "none";
defparam ram_block1a29.port_a_data_out_clock = "none";
defparam ram_block1a29.port_a_data_width = 1;
defparam ram_block1a29.port_a_first_address = 0;
defparam ram_block1a29.port_a_first_bit_number = 29;
defparam ram_block1a29.port_a_last_address = 1023;
defparam ram_block1a29.port_a_logical_ram_depth = 1024;
defparam ram_block1a29.port_a_logical_ram_width = 32;
defparam ram_block1a29.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a29.ram_block_type = "auto";
defparam ram_block1a29.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a13(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a13_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a13.init_file_layout = "port_a";
defparam ram_block1a13.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.operation_mode = "single_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 10;
defparam ram_block1a13.port_a_byte_enable_mask_width = 1;
defparam ram_block1a13.port_a_byte_size = 1;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 1023;
defparam ram_block1a13.port_a_logical_ram_depth = 1024;
defparam ram_block1a13.port_a_logical_ram_width = 32;
defparam ram_block1a13.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a13.ram_block_type = "auto";
defparam ram_block1a13.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a28(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[28]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a28_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a28.clk0_core_clock_enable = "ena0";
defparam ram_block1a28.clk0_input_clock_enable = "ena0";
defparam ram_block1a28.data_interleave_offset_in_bits = 1;
defparam ram_block1a28.data_interleave_width_in_bits = 1;
defparam ram_block1a28.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a28.init_file_layout = "port_a";
defparam ram_block1a28.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a28.operation_mode = "single_port";
defparam ram_block1a28.port_a_address_clear = "none";
defparam ram_block1a28.port_a_address_width = 10;
defparam ram_block1a28.port_a_byte_enable_mask_width = 1;
defparam ram_block1a28.port_a_byte_size = 1;
defparam ram_block1a28.port_a_data_out_clear = "none";
defparam ram_block1a28.port_a_data_out_clock = "none";
defparam ram_block1a28.port_a_data_width = 1;
defparam ram_block1a28.port_a_first_address = 0;
defparam ram_block1a28.port_a_first_bit_number = 28;
defparam ram_block1a28.port_a_last_address = 1023;
defparam ram_block1a28.port_a_logical_ram_depth = 1024;
defparam ram_block1a28.port_a_logical_ram_width = 32;
defparam ram_block1a28.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a28.ram_block_type = "auto";
defparam ram_block1a28.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a12(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a12_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a12.init_file_layout = "port_a";
defparam ram_block1a12.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.operation_mode = "single_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 10;
defparam ram_block1a12.port_a_byte_enable_mask_width = 1;
defparam ram_block1a12.port_a_byte_size = 1;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 1023;
defparam ram_block1a12.port_a_logical_ram_depth = 1024;
defparam ram_block1a12.port_a_logical_ram_width = 32;
defparam ram_block1a12.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a12.ram_block_type = "auto";
defparam ram_block1a12.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a27(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[27]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a27_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a27.clk0_core_clock_enable = "ena0";
defparam ram_block1a27.clk0_input_clock_enable = "ena0";
defparam ram_block1a27.data_interleave_offset_in_bits = 1;
defparam ram_block1a27.data_interleave_width_in_bits = 1;
defparam ram_block1a27.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a27.init_file_layout = "port_a";
defparam ram_block1a27.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a27.operation_mode = "single_port";
defparam ram_block1a27.port_a_address_clear = "none";
defparam ram_block1a27.port_a_address_width = 10;
defparam ram_block1a27.port_a_byte_enable_mask_width = 1;
defparam ram_block1a27.port_a_byte_size = 1;
defparam ram_block1a27.port_a_data_out_clear = "none";
defparam ram_block1a27.port_a_data_out_clock = "none";
defparam ram_block1a27.port_a_data_width = 1;
defparam ram_block1a27.port_a_first_address = 0;
defparam ram_block1a27.port_a_first_bit_number = 27;
defparam ram_block1a27.port_a_last_address = 1023;
defparam ram_block1a27.port_a_logical_ram_depth = 1024;
defparam ram_block1a27.port_a_logical_ram_width = 32;
defparam ram_block1a27.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a27.ram_block_type = "auto";
defparam ram_block1a27.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a11(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a11_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a11.init_file_layout = "port_a";
defparam ram_block1a11.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.operation_mode = "single_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 10;
defparam ram_block1a11.port_a_byte_enable_mask_width = 1;
defparam ram_block1a11.port_a_byte_size = 1;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 1023;
defparam ram_block1a11.port_a_logical_ram_depth = 1024;
defparam ram_block1a11.port_a_logical_ram_width = 32;
defparam ram_block1a11.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a11.ram_block_type = "auto";
defparam ram_block1a11.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a25(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[25]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a25_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a25.clk0_core_clock_enable = "ena0";
defparam ram_block1a25.clk0_input_clock_enable = "ena0";
defparam ram_block1a25.data_interleave_offset_in_bits = 1;
defparam ram_block1a25.data_interleave_width_in_bits = 1;
defparam ram_block1a25.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a25.init_file_layout = "port_a";
defparam ram_block1a25.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a25.operation_mode = "single_port";
defparam ram_block1a25.port_a_address_clear = "none";
defparam ram_block1a25.port_a_address_width = 10;
defparam ram_block1a25.port_a_byte_enable_mask_width = 1;
defparam ram_block1a25.port_a_byte_size = 1;
defparam ram_block1a25.port_a_data_out_clear = "none";
defparam ram_block1a25.port_a_data_out_clock = "none";
defparam ram_block1a25.port_a_data_width = 1;
defparam ram_block1a25.port_a_first_address = 0;
defparam ram_block1a25.port_a_first_bit_number = 25;
defparam ram_block1a25.port_a_last_address = 1023;
defparam ram_block1a25.port_a_logical_ram_depth = 1024;
defparam ram_block1a25.port_a_logical_ram_width = 32;
defparam ram_block1a25.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a25.ram_block_type = "auto";
defparam ram_block1a25.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a9(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a9_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a9.init_file_layout = "port_a";
defparam ram_block1a9.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.operation_mode = "single_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 10;
defparam ram_block1a9.port_a_byte_enable_mask_width = 1;
defparam ram_block1a9.port_a_byte_size = 1;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 1023;
defparam ram_block1a9.port_a_logical_ram_depth = 1024;
defparam ram_block1a9.port_a_logical_ram_width = 32;
defparam ram_block1a9.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a9.ram_block_type = "auto";
defparam ram_block1a9.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a24(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[24]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a24_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a24.clk0_core_clock_enable = "ena0";
defparam ram_block1a24.clk0_input_clock_enable = "ena0";
defparam ram_block1a24.data_interleave_offset_in_bits = 1;
defparam ram_block1a24.data_interleave_width_in_bits = 1;
defparam ram_block1a24.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a24.init_file_layout = "port_a";
defparam ram_block1a24.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a24.operation_mode = "single_port";
defparam ram_block1a24.port_a_address_clear = "none";
defparam ram_block1a24.port_a_address_width = 10;
defparam ram_block1a24.port_a_byte_enable_mask_width = 1;
defparam ram_block1a24.port_a_byte_size = 1;
defparam ram_block1a24.port_a_data_out_clear = "none";
defparam ram_block1a24.port_a_data_out_clock = "none";
defparam ram_block1a24.port_a_data_width = 1;
defparam ram_block1a24.port_a_first_address = 0;
defparam ram_block1a24.port_a_first_bit_number = 24;
defparam ram_block1a24.port_a_last_address = 1023;
defparam ram_block1a24.port_a_logical_ram_depth = 1024;
defparam ram_block1a24.port_a_logical_ram_width = 32;
defparam ram_block1a24.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a24.ram_block_type = "auto";
defparam ram_block1a24.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a8(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a8_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a8.init_file_layout = "port_a";
defparam ram_block1a8.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.operation_mode = "single_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 10;
defparam ram_block1a8.port_a_byte_enable_mask_width = 1;
defparam ram_block1a8.port_a_byte_size = 1;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 1023;
defparam ram_block1a8.port_a_logical_ram_depth = 1024;
defparam ram_block1a8.port_a_logical_ram_width = 32;
defparam ram_block1a8.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a8.ram_block_type = "auto";
defparam ram_block1a8.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a6(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.operation_mode = "single_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 10;
defparam ram_block1a6.port_a_byte_enable_mask_width = 1;
defparam ram_block1a6.port_a_byte_size = 1;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 1023;
defparam ram_block1a6.port_a_logical_ram_depth = 1024;
defparam ram_block1a6.port_a_logical_ram_width = 32;
defparam ram_block1a6.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a14(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[1]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a14_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a14.init_file_layout = "port_a";
defparam ram_block1a14.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.operation_mode = "single_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 10;
defparam ram_block1a14.port_a_byte_enable_mask_width = 1;
defparam ram_block1a14.port_a_byte_size = 1;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 1023;
defparam ram_block1a14.port_a_logical_ram_depth = 1024;
defparam ram_block1a14.port_a_logical_ram_width = 32;
defparam ram_block1a14.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a14.ram_block_type = "auto";
defparam ram_block1a14.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a22(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[22]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a22_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a22.clk0_core_clock_enable = "ena0";
defparam ram_block1a22.clk0_input_clock_enable = "ena0";
defparam ram_block1a22.data_interleave_offset_in_bits = 1;
defparam ram_block1a22.data_interleave_width_in_bits = 1;
defparam ram_block1a22.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a22.init_file_layout = "port_a";
defparam ram_block1a22.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a22.operation_mode = "single_port";
defparam ram_block1a22.port_a_address_clear = "none";
defparam ram_block1a22.port_a_address_width = 10;
defparam ram_block1a22.port_a_byte_enable_mask_width = 1;
defparam ram_block1a22.port_a_byte_size = 1;
defparam ram_block1a22.port_a_data_out_clear = "none";
defparam ram_block1a22.port_a_data_out_clock = "none";
defparam ram_block1a22.port_a_data_width = 1;
defparam ram_block1a22.port_a_first_address = 0;
defparam ram_block1a22.port_a_first_bit_number = 22;
defparam ram_block1a22.port_a_last_address = 1023;
defparam ram_block1a22.port_a_logical_ram_depth = 1024;
defparam ram_block1a22.port_a_logical_ram_width = 32;
defparam ram_block1a22.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a22.ram_block_type = "auto";
defparam ram_block1a22.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a30(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[30]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[3]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a30_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a30.clk0_core_clock_enable = "ena0";
defparam ram_block1a30.clk0_input_clock_enable = "ena0";
defparam ram_block1a30.data_interleave_offset_in_bits = 1;
defparam ram_block1a30.data_interleave_width_in_bits = 1;
defparam ram_block1a30.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a30.init_file_layout = "port_a";
defparam ram_block1a30.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a30.operation_mode = "single_port";
defparam ram_block1a30.port_a_address_clear = "none";
defparam ram_block1a30.port_a_address_width = 10;
defparam ram_block1a30.port_a_byte_enable_mask_width = 1;
defparam ram_block1a30.port_a_byte_size = 1;
defparam ram_block1a30.port_a_data_out_clear = "none";
defparam ram_block1a30.port_a_data_out_clock = "none";
defparam ram_block1a30.port_a_data_width = 1;
defparam ram_block1a30.port_a_first_address = 0;
defparam ram_block1a30.port_a_first_bit_number = 30;
defparam ram_block1a30.port_a_last_address = 1023;
defparam ram_block1a30.port_a_logical_ram_depth = 1024;
defparam ram_block1a30.port_a_logical_ram_width = 32;
defparam ram_block1a30.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a30.ram_block_type = "auto";
defparam ram_block1a30.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a5(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.operation_mode = "single_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 10;
defparam ram_block1a5.port_a_byte_enable_mask_width = 1;
defparam ram_block1a5.port_a_byte_size = 1;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 1023;
defparam ram_block1a5.port_a_logical_ram_depth = 1024;
defparam ram_block1a5.port_a_logical_ram_width = 32;
defparam ram_block1a5.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a21(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[21]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a21_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a21.clk0_core_clock_enable = "ena0";
defparam ram_block1a21.clk0_input_clock_enable = "ena0";
defparam ram_block1a21.data_interleave_offset_in_bits = 1;
defparam ram_block1a21.data_interleave_width_in_bits = 1;
defparam ram_block1a21.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a21.init_file_layout = "port_a";
defparam ram_block1a21.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a21.operation_mode = "single_port";
defparam ram_block1a21.port_a_address_clear = "none";
defparam ram_block1a21.port_a_address_width = 10;
defparam ram_block1a21.port_a_byte_enable_mask_width = 1;
defparam ram_block1a21.port_a_byte_size = 1;
defparam ram_block1a21.port_a_data_out_clear = "none";
defparam ram_block1a21.port_a_data_out_clock = "none";
defparam ram_block1a21.port_a_data_width = 1;
defparam ram_block1a21.port_a_first_address = 0;
defparam ram_block1a21.port_a_first_bit_number = 21;
defparam ram_block1a21.port_a_last_address = 1023;
defparam ram_block1a21.port_a_logical_ram_depth = 1024;
defparam ram_block1a21.port_a_logical_ram_width = 32;
defparam ram_block1a21.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a21.ram_block_type = "auto";
defparam ram_block1a21.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a4(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.operation_mode = "single_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 10;
defparam ram_block1a4.port_a_byte_enable_mask_width = 1;
defparam ram_block1a4.port_a_byte_size = 1;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 1023;
defparam ram_block1a4.port_a_logical_ram_depth = 1024;
defparam ram_block1a4.port_a_logical_ram_width = 32;
defparam ram_block1a4.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a20(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[20]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a20_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a20.clk0_core_clock_enable = "ena0";
defparam ram_block1a20.clk0_input_clock_enable = "ena0";
defparam ram_block1a20.data_interleave_offset_in_bits = 1;
defparam ram_block1a20.data_interleave_width_in_bits = 1;
defparam ram_block1a20.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a20.init_file_layout = "port_a";
defparam ram_block1a20.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a20.operation_mode = "single_port";
defparam ram_block1a20.port_a_address_clear = "none";
defparam ram_block1a20.port_a_address_width = 10;
defparam ram_block1a20.port_a_byte_enable_mask_width = 1;
defparam ram_block1a20.port_a_byte_size = 1;
defparam ram_block1a20.port_a_data_out_clear = "none";
defparam ram_block1a20.port_a_data_out_clock = "none";
defparam ram_block1a20.port_a_data_width = 1;
defparam ram_block1a20.port_a_first_address = 0;
defparam ram_block1a20.port_a_first_bit_number = 20;
defparam ram_block1a20.port_a_last_address = 1023;
defparam ram_block1a20.port_a_logical_ram_depth = 1024;
defparam ram_block1a20.port_a_logical_ram_width = 32;
defparam ram_block1a20.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a20.ram_block_type = "auto";
defparam ram_block1a20.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a3(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.operation_mode = "single_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 10;
defparam ram_block1a3.port_a_byte_enable_mask_width = 1;
defparam ram_block1a3.port_a_byte_size = 1;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 1023;
defparam ram_block1a3.port_a_logical_ram_depth = 1024;
defparam ram_block1a3.port_a_logical_ram_width = 32;
defparam ram_block1a3.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a19(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[19]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a19_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a19.clk0_core_clock_enable = "ena0";
defparam ram_block1a19.clk0_input_clock_enable = "ena0";
defparam ram_block1a19.data_interleave_offset_in_bits = 1;
defparam ram_block1a19.data_interleave_width_in_bits = 1;
defparam ram_block1a19.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a19.init_file_layout = "port_a";
defparam ram_block1a19.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a19.operation_mode = "single_port";
defparam ram_block1a19.port_a_address_clear = "none";
defparam ram_block1a19.port_a_address_width = 10;
defparam ram_block1a19.port_a_byte_enable_mask_width = 1;
defparam ram_block1a19.port_a_byte_size = 1;
defparam ram_block1a19.port_a_data_out_clear = "none";
defparam ram_block1a19.port_a_data_out_clock = "none";
defparam ram_block1a19.port_a_data_width = 1;
defparam ram_block1a19.port_a_first_address = 0;
defparam ram_block1a19.port_a_first_bit_number = 19;
defparam ram_block1a19.port_a_last_address = 1023;
defparam ram_block1a19.port_a_logical_ram_depth = 1024;
defparam ram_block1a19.port_a_logical_ram_width = 32;
defparam ram_block1a19.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a19.ram_block_type = "auto";
defparam ram_block1a19.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a1(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.operation_mode = "single_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 10;
defparam ram_block1a1.port_a_byte_enable_mask_width = 1;
defparam ram_block1a1.port_a_byte_size = 1;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 1023;
defparam ram_block1a1.port_a_logical_ram_depth = 1024;
defparam ram_block1a1.port_a_logical_ram_width = 32;
defparam ram_block1a1.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a17(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[17]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a17_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a17.clk0_core_clock_enable = "ena0";
defparam ram_block1a17.clk0_input_clock_enable = "ena0";
defparam ram_block1a17.data_interleave_offset_in_bits = 1;
defparam ram_block1a17.data_interleave_width_in_bits = 1;
defparam ram_block1a17.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a17.init_file_layout = "port_a";
defparam ram_block1a17.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a17.operation_mode = "single_port";
defparam ram_block1a17.port_a_address_clear = "none";
defparam ram_block1a17.port_a_address_width = 10;
defparam ram_block1a17.port_a_byte_enable_mask_width = 1;
defparam ram_block1a17.port_a_byte_size = 1;
defparam ram_block1a17.port_a_data_out_clear = "none";
defparam ram_block1a17.port_a_data_out_clock = "none";
defparam ram_block1a17.port_a_data_width = 1;
defparam ram_block1a17.port_a_first_address = 0;
defparam ram_block1a17.port_a_first_bit_number = 17;
defparam ram_block1a17.port_a_last_address = 1023;
defparam ram_block1a17.port_a_logical_ram_depth = 1024;
defparam ram_block1a17.port_a_logical_ram_width = 32;
defparam ram_block1a17.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a17.ram_block_type = "auto";
defparam ram_block1a17.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a0(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[0]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.operation_mode = "single_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 10;
defparam ram_block1a0.port_a_byte_enable_mask_width = 1;
defparam ram_block1a0.port_a_byte_size = 1;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 1023;
defparam ram_block1a0.port_a_logical_ram_depth = 1024;
defparam ram_block1a0.port_a_logical_ram_width = 32;
defparam ram_block1a0.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

cyclonev_ram_block ram_block1a16(
	.portawe(!wren_a),
	.portare(wren_a),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(!clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.nerror(vcc),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[16]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,byteena_a[2]}),
	.portbdatain(1'b0),
	.portbaddr(1'b0),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a16_PORTADATAOUT_bus),
	.portbdataout(),
	.eccstatus(),
	.dftout());
defparam ram_block1a16.clk0_core_clock_enable = "ena0";
defparam ram_block1a16.clk0_input_clock_enable = "ena0";
defparam ram_block1a16.data_interleave_offset_in_bits = 1;
defparam ram_block1a16.data_interleave_width_in_bits = 1;
defparam ram_block1a16.init_file = "embedded_system_onchip_memory2_0.hex";
defparam ram_block1a16.init_file_layout = "port_a";
defparam ram_block1a16.logical_ram_name = "embedded_system_onchip_memory2_0:onchip_memory2_0|altsyncram:the_altsyncram|altsyncram_45o1:auto_generated|ALTSYNCRAM";
defparam ram_block1a16.operation_mode = "single_port";
defparam ram_block1a16.port_a_address_clear = "none";
defparam ram_block1a16.port_a_address_width = 10;
defparam ram_block1a16.port_a_byte_enable_mask_width = 1;
defparam ram_block1a16.port_a_byte_size = 1;
defparam ram_block1a16.port_a_data_out_clear = "none";
defparam ram_block1a16.port_a_data_out_clock = "none";
defparam ram_block1a16.port_a_data_width = 1;
defparam ram_block1a16.port_a_first_address = 0;
defparam ram_block1a16.port_a_first_bit_number = 16;
defparam ram_block1a16.port_a_last_address = 1023;
defparam ram_block1a16.port_a_logical_ram_depth = 1024;
defparam ram_block1a16.port_a_logical_ram_width = 32;
defparam ram_block1a16.port_a_read_during_write_mode = "dont_care";
defparam ram_block1a16.ram_block_type = "auto";
defparam ram_block1a16.mem_init0 = "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";

endmodule
