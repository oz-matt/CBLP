
module embedded_system (
	clk_clk,
	ad9833_io_readdata);	

	input		clk_clk;
	output	[31:0]	ad9833_io_readdata;
endmodule
